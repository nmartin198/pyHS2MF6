time,SOUTHOUT
1.000000000000,-202.28
2.000000000000,-202.44
3.000000000000,-201.91
4.000000000000,-201.44
5.000000000000,-200.30
6.000000000000,-198.87
7.000000000000,-197.62
8.000000000000,-196.50
9.000000000000,-198.42
10.00000000000,-198.90
11.00000000000,-195.09
12.00000000000,-193.48
13.00000000000,-192.32
14.00000000000,-191.37
15.00000000000,-190.48
16.00000000000,-189.66
17.00000000000,-188.89
18.00000000000,-188.17
19.00000000000,-187.47
20.00000000000,-186.81
21.00000000000,-186.18
22.00000000000,-185.58
23.00000000000,-185.00
24.00000000000,-184.46
25.00000000000,-183.93
26.00000000000,-183.42
27.00000000000,-182.93
28.00000000000,-182.45
29.00000000000,-181.98
30.00000000000,-181.53
31.00000000000,-181.08
32.00000000000,-180.65
33.00000000000,-180.22
34.00000000000,-179.81
35.00000000000,-179.41
36.00000000000,-179.01
37.00000000000,-178.62
38.00000000000,-178.25
39.00000000000,-177.88
40.00000000000,-177.51
41.00000000000,-177.17
42.00000000000,-176.82
43.00000000000,-176.48
44.00000000000,-176.14
45.00000000000,-175.81
46.00000000000,-175.49
47.00000000000,-175.17
48.00000000000,-174.87
49.00000000000,-174.58
50.00000000000,-174.29
51.00000000000,-174.01
52.00000000000,-173.76
53.00000000000,-173.47
54.00000000000,-173.19
55.00000000000,-172.92
56.00000000000,-172.68
57.00000000000,-172.41
58.00000000000,-172.14
59.00000000000,-171.87
60.00000000000,-171.62
61.00000000000,-171.37
62.00000000000,-171.12
63.00000000000,-170.88
64.00000000000,-170.64
65.00000000000,-170.40
66.00000000000,-170.16
67.00000000000,-169.92
68.00000000000,-169.69
69.00000000000,-169.55
70.00000000000,-169.29
71.00000000000,-169.04
72.00000000000,-168.81
73.00000000000,-168.58
74.00000000000,-168.36
75.00000000000,-168.14
76.00000000000,-167.93
77.00000000000,-167.72
78.00000000000,-167.51
79.00000000000,-167.30
80.00000000000,-167.09
81.00000000000,-166.89
82.00000000000,-166.72
83.00000000000,-166.51
84.00000000000,-166.29
85.00000000000,-166.09
86.00000000000,-165.89
87.00000000000,-165.69
88.00000000000,-165.49
89.00000000000,-165.30
90.00000000000,-165.11
91.00000000000,-164.91
92.00000000000,-164.72
93.00000000000,-164.70
94.00000000000,-164.45
95.00000000000,-164.22
96.00000000000,-164.00
97.00000000000,-163.79
98.00000000000,-163.59
99.00000000000,-163.39
100.0000000000,-163.20
101.0000000000,-163.01
102.0000000000,-162.82
103.0000000000,-162.63
104.0000000000,-162.44
105.0000000000,-162.25
106.0000000000,-162.06
107.0000000000,-161.88
108.0000000000,-161.78
109.0000000000,-161.57
110.0000000000,-161.36
111.0000000000,-161.17
112.0000000000,-160.98
113.0000000000,-160.80
114.0000000000,-160.62
115.0000000000,-160.45
116.0000000000,-160.27
117.0000000000,-160.10
118.0000000000,-160.19
119.0000000000,-160.39
120.0000000000,-159.97
121.0000000000,-159.63
122.0000000000,-159.55
123.0000000000,-159.27
124.0000000000,-159.04
125.0000000000,-158.84
126.0000000000,-158.66
127.0000000000,-158.49
128.0000000000,-158.32
129.0000000000,-158.15
130.0000000000,-158.06
131.0000000000,-157.96
132.0000000000,-157.74
133.0000000000,-157.55
134.0000000000,-157.37
135.0000000000,-157.32
136.0000000000,-157.11
137.0000000000,-156.92
138.0000000000,-156.75
139.0000000000,-156.58
140.0000000000,-156.42
141.0000000000,-156.27
142.0000000000,-156.11
143.0000000000,-155.95
144.0000000000,-156.04
145.0000000000,-155.81
146.0000000000,-156.02
147.0000000000,-155.66
148.0000000000,-155.39
149.0000000000,-155.22
150.0000000000,-155.02
151.0000000000,-154.84
152.0000000000,-154.68
153.0000000000,-154.53
154.0000000000,-154.38
155.0000000000,-154.23
156.0000000000,-154.08
157.0000000000,-153.94
158.0000000000,-153.79
159.0000000000,-153.72
160.0000000000,-153.55
161.0000000000,-153.39
162.0000000000,-153.23
163.0000000000,-153.09
164.0000000000,-152.94
165.0000000000,-152.85
166.0000000000,-153.13
167.0000000000,-152.84
168.0000000000,-152.57
169.0000000000,-152.40
170.0000000000,-152.22
171.0000000000,-152.06
172.0000000000,-151.91
173.0000000000,-151.77
174.0000000000,-151.63
175.0000000000,-151.49
176.0000000000,-151.36
177.0000000000,-151.22
178.0000000000,-151.09
179.0000000000,-150.95
180.0000000000,-150.82
181.0000000000,-150.76
182.0000000000,-150.60
183.0000000000,-150.47
184.0000000000,-150.32
185.0000000000,-150.19
186.0000000000,-150.05
187.0000000000,-149.92
188.0000000000,-149.79
189.0000000000,-149.66
190.0000000000,-149.53
191.0000000000,-149.41
192.0000000000,-149.28
193.0000000000,-149.15
194.0000000000,-149.03
195.0000000000,-148.90
196.0000000000,-148.79
197.0000000000,-148.84
198.0000000000,-148.73
199.0000000000,-148.55
200.0000000000,-148.41
201.0000000000,-148.25
202.0000000000,-148.11
203.0000000000,-147.99
204.0000000000,-147.86
205.0000000000,-147.73
206.0000000000,-147.61
207.0000000000,-147.49
208.0000000000,-147.37
209.0000000000,-147.25
210.0000000000,-147.15
211.0000000000,-147.02
212.0000000000,-146.90
213.0000000000,-146.78
214.0000000000,-146.66
215.0000000000,-146.54
216.0000000000,-146.43
217.0000000000,-146.31
218.0000000000,-146.19
219.0000000000,-146.08
220.0000000000,-145.96
221.0000000000,-145.85
222.0000000000,-145.73
223.0000000000,-145.62
224.0000000000,-145.51
225.0000000000,-145.39
226.0000000000,-145.28
227.0000000000,-145.16
228.0000000000,-145.05
229.0000000000,-144.94
230.0000000000,-144.83
231.0000000000,-144.71
232.0000000000,-144.60
233.0000000000,-144.49
234.0000000000,-144.38
235.0000000000,-144.27
236.0000000000,-144.27
237.0000000000,-144.12
238.0000000000,-144.00
239.0000000000,-144.02
240.0000000000,-143.96
241.0000000000,-143.77
242.0000000000,-143.63
243.0000000000,-143.50
244.0000000000,-143.39
245.0000000000,-143.28
246.0000000000,-143.22
247.0000000000,-143.09
248.0000000000,-143.01
249.0000000000,-142.91
250.0000000000,-142.78
251.0000000000,-142.67
252.0000000000,-142.59
253.0000000000,-142.47
254.0000000000,-142.37
255.0000000000,-142.26
256.0000000000,-142.15
257.0000000000,-142.04
258.0000000000,-141.94
259.0000000000,-141.84
260.0000000000,-141.76
261.0000000000,-141.69
262.0000000000,-141.58
263.0000000000,-141.77
264.0000000000,-141.78
265.0000000000,-141.51
266.0000000000,-141.33
267.0000000000,-141.20
268.0000000000,-141.09
269.0000000000,-140.98
270.0000000000,-140.87
271.0000000000,-140.77
272.0000000000,-140.70
273.0000000000,-140.59
274.0000000000,-140.49
275.0000000000,-140.39
276.0000000000,-140.29
277.0000000000,-140.19
278.0000000000,-140.09
279.0000000000,-139.99
280.0000000000,-139.89
281.0000000000,-139.80
282.0000000000,-139.70
283.0000000000,-139.60
284.0000000000,-139.51
285.0000000000,-139.41
286.0000000000,-139.32
287.0000000000,-139.23
288.0000000000,-139.16
289.0000000000,-139.22
290.0000000000,-139.06
291.0000000000,-138.94
292.0000000000,-138.83
293.0000000000,-138.73
294.0000000000,-138.63
295.0000000000,-138.53
296.0000000000,-138.44
297.0000000000,-138.35
298.0000000000,-138.25
299.0000000000,-138.16
300.0000000000,-138.07
301.0000000000,-137.98
302.0000000000,-137.88
303.0000000000,-137.79
304.0000000000,-137.70
305.0000000000,-137.61
306.0000000000,-137.52
307.0000000000,-137.43
308.0000000000,-137.34
309.0000000000,-137.25
310.0000000000,-137.17
311.0000000000,-137.08
312.0000000000,-137.00
313.0000000000,-136.91
314.0000000000,-136.82
315.0000000000,-136.73
316.0000000000,-136.64
317.0000000000,-136.55
318.0000000000,-136.47
319.0000000000,-136.38
320.0000000000,-136.29
321.0000000000,-136.20
322.0000000000,-136.11
323.0000000000,-136.03
324.0000000000,-135.94
325.0000000000,-135.85
326.0000000000,-135.77
327.0000000000,-135.68
328.0000000000,-135.61
329.0000000000,-135.53
330.0000000000,-135.45
331.0000000000,-135.36
332.0000000000,-135.28
333.0000000000,-135.19
334.0000000000,-135.10
335.0000000000,-135.02
336.0000000000,-134.93
337.0000000000,-134.85
338.0000000000,-134.77
339.0000000000,-134.68
340.0000000000,-134.60
341.0000000000,-134.52
342.0000000000,-134.43
343.0000000000,-134.35
344.0000000000,-134.27
345.0000000000,-134.18
346.0000000000,-134.10
347.0000000000,-134.02
348.0000000000,-133.93
349.0000000000,-133.85
350.0000000000,-133.77
351.0000000000,-133.69
352.0000000000,-133.61
353.0000000000,-133.52
354.0000000000,-133.44
355.0000000000,-133.37
356.0000000000,-133.29
357.0000000000,-133.21
358.0000000000,-133.13
359.0000000000,-133.05
360.0000000000,-132.97
361.0000000000,-132.90
362.0000000000,-132.82
363.0000000000,-132.74
364.0000000000,-132.66
365.0000000000,-132.58
366.0000000000,-132.50
367.0000000000,-132.43
368.0000000000,-132.35
369.0000000000,-132.27
370.0000000000,-132.19
371.0000000000,-132.11
372.0000000000,-132.03
373.0000000000,-131.95
374.0000000000,-131.88
375.0000000000,-131.80
376.0000000000,-131.72
377.0000000000,-131.64
378.0000000000,-131.57
379.0000000000,-131.49
380.0000000000,-131.41
381.0000000000,-131.33
382.0000000000,-131.26
383.0000000000,-131.18
384.0000000000,-131.11
385.0000000000,-131.03
386.0000000000,-130.95
387.0000000000,-130.88
388.0000000000,-130.80
389.0000000000,-130.73
390.0000000000,-130.65
391.0000000000,-130.58
392.0000000000,-130.50
393.0000000000,-130.43
394.0000000000,-130.35
395.0000000000,-130.28
396.0000000000,-130.20
397.0000000000,-130.13
398.0000000000,-130.05
399.0000000000,-129.98
400.0000000000,-129.90
401.0000000000,-129.83
402.0000000000,-129.76
403.0000000000,-129.68
404.0000000000,-129.61
405.0000000000,-129.54
406.0000000000,-129.46
407.0000000000,-129.39
408.0000000000,-129.32
409.0000000000,-129.24
410.0000000000,-129.17
411.0000000000,-129.10
412.0000000000,-129.03
413.0000000000,-128.96
414.0000000000,-128.88
415.0000000000,-128.81
416.0000000000,-128.74
417.0000000000,-128.67
418.0000000000,-128.60
419.0000000000,-128.53
420.0000000000,-128.45
421.0000000000,-128.38
422.0000000000,-128.32
423.0000000000,-128.25
424.0000000000,-128.18
425.0000000000,-128.11
426.0000000000,-128.04
427.0000000000,-127.97
428.0000000000,-127.90
429.0000000000,-127.83
430.0000000000,-127.76
431.0000000000,-127.69
432.0000000000,-127.62
433.0000000000,-127.55
434.0000000000,-127.48
435.0000000000,-127.41
436.0000000000,-127.34
437.0000000000,-127.27
438.0000000000,-127.21
439.0000000000,-127.14
440.0000000000,-127.07
441.0000000000,-127.00
442.0000000000,-126.93
443.0000000000,-126.86
444.0000000000,-126.79
445.0000000000,-126.73
446.0000000000,-126.66
447.0000000000,-126.59
448.0000000000,-126.52
449.0000000000,-126.46
450.0000000000,-126.39
451.0000000000,-126.32
452.0000000000,-126.26
453.0000000000,-126.19
454.0000000000,-126.12
455.0000000000,-126.06
456.0000000000,-125.99
457.0000000000,-125.92
458.0000000000,-125.86
459.0000000000,-125.79
460.0000000000,-125.73
461.0000000000,-125.66
462.0000000000,-125.60
463.0000000000,-125.53
464.0000000000,-125.47
465.0000000000,-125.40
466.0000000000,-125.34
467.0000000000,-125.27
468.0000000000,-125.20
469.0000000000,-125.14
470.0000000000,-125.07
471.0000000000,-125.01
472.0000000000,-124.94
473.0000000000,-124.88
474.0000000000,-124.82
475.0000000000,-124.75
476.0000000000,-124.69
477.0000000000,-124.62
478.0000000000,-124.56
479.0000000000,-124.49
480.0000000000,-124.43
481.0000000000,-124.37
482.0000000000,-124.30
483.0000000000,-124.24
484.0000000000,-124.18
485.0000000000,-124.11
486.0000000000,-124.05
487.0000000000,-123.99
488.0000000000,-123.92
489.0000000000,-123.86
490.0000000000,-123.80
491.0000000000,-123.73
492.0000000000,-123.68
493.0000000000,-123.61
494.0000000000,-123.55
495.0000000000,-123.49
496.0000000000,-123.43
497.0000000000,-123.37
498.0000000000,-123.31
499.0000000000,-123.25
500.0000000000,-123.19
501.0000000000,-123.13
502.0000000000,-123.07
503.0000000000,-123.01
504.0000000000,-122.94
505.0000000000,-122.88
506.0000000000,-122.82
507.0000000000,-122.76
508.0000000000,-122.70
509.0000000000,-122.64
510.0000000000,-122.58
511.0000000000,-122.54
512.0000000000,-122.49
513.0000000000,-122.43
514.0000000000,-122.37
515.0000000000,-122.31
516.0000000000,-122.25
517.0000000000,-122.19
518.0000000000,-122.13
519.0000000000,-122.07
520.0000000000,-122.01
521.0000000000,-121.95
522.0000000000,-121.89
523.0000000000,-121.83
524.0000000000,-121.77
525.0000000000,-121.71
526.0000000000,-121.65
527.0000000000,-121.59
528.0000000000,-121.53
529.0000000000,-121.48
530.0000000000,-121.43
531.0000000000,-121.37
532.0000000000,-121.32
533.0000000000,-121.26
534.0000000000,-121.20
535.0000000000,-121.14
536.0000000000,-121.13
537.0000000000,-121.10
538.0000000000,-121.05
539.0000000000,-121.00
540.0000000000,-120.94
541.0000000000,-120.90
542.0000000000,-120.85
543.0000000000,-120.79
544.0000000000,-120.73
545.0000000000,-120.68
546.0000000000,-120.62
547.0000000000,-120.56
548.0000000000,-120.50
549.0000000000,-120.45
550.0000000000,-120.39
551.0000000000,-120.33
552.0000000000,-120.27
553.0000000000,-120.22
554.0000000000,-120.16
555.0000000000,-120.10
556.0000000000,-120.05
557.0000000000,-119.99
558.0000000000,-119.94
559.0000000000,-119.88
560.0000000000,-119.83
561.0000000000,-119.77
562.0000000000,-119.72
563.0000000000,-119.67
564.0000000000,-119.62
565.0000000000,-119.56
566.0000000000,-119.51
567.0000000000,-119.45
568.0000000000,-119.40
569.0000000000,-119.34
570.0000000000,-119.28
571.0000000000,-119.23
572.0000000000,-119.18
573.0000000000,-119.12
574.0000000000,-119.06
575.0000000000,-119.01
576.0000000000,-118.95
577.0000000000,-118.90
578.0000000000,-118.84
579.0000000000,-118.80
580.0000000000,-118.77
581.0000000000,-118.72
582.0000000000,-118.66
583.0000000000,-118.61
584.0000000000,-118.56
585.0000000000,-118.50
586.0000000000,-118.45
587.0000000000,-118.39
588.0000000000,-118.34
589.0000000000,-118.29
590.0000000000,-118.24
591.0000000000,-118.19
592.0000000000,-118.13
593.0000000000,-118.08
594.0000000000,-118.03
595.0000000000,-117.98
596.0000000000,-117.93
597.0000000000,-117.88
598.0000000000,-117.83
599.0000000000,-117.78
600.0000000000,-117.73
601.0000000000,-117.67
602.0000000000,-117.62
603.0000000000,-117.57
604.0000000000,-117.51
605.0000000000,-117.46
606.0000000000,-117.41
607.0000000000,-117.36
608.0000000000,-117.30
609.0000000000,-117.25
610.0000000000,-117.20
611.0000000000,-117.15
612.0000000000,-117.09
613.0000000000,-117.05
614.0000000000,-117.00
615.0000000000,-116.95
616.0000000000,-116.90
617.0000000000,-116.85
618.0000000000,-116.80
619.0000000000,-116.75
620.0000000000,-116.70
621.0000000000,-116.65
622.0000000000,-116.60
623.0000000000,-116.55
624.0000000000,-116.50
625.0000000000,-116.45
626.0000000000,-116.39
627.0000000000,-116.35
628.0000000000,-116.31
629.0000000000,-116.26
630.0000000000,-116.22
631.0000000000,-116.17
632.0000000000,-116.12
633.0000000000,-116.07
634.0000000000,-116.02
635.0000000000,-115.99
636.0000000000,-115.95
637.0000000000,-115.90
638.0000000000,-115.85
639.0000000000,-115.80
640.0000000000,-115.75
641.0000000000,-115.70
642.0000000000,-115.65
643.0000000000,-115.60
644.0000000000,-115.55
645.0000000000,-115.50
646.0000000000,-115.45
647.0000000000,-115.40
648.0000000000,-115.35
649.0000000000,-115.31
650.0000000000,-115.26
651.0000000000,-115.22
652.0000000000,-115.17
653.0000000000,-115.12
654.0000000000,-115.07
655.0000000000,-115.02
656.0000000000,-114.97
657.0000000000,-114.92
658.0000000000,-114.87
659.0000000000,-114.82
660.0000000000,-114.78
661.0000000000,-114.73
662.0000000000,-114.69
663.0000000000,-114.64
664.0000000000,-114.59
665.0000000000,-114.54
666.0000000000,-114.49
667.0000000000,-114.44
668.0000000000,-114.40
669.0000000000,-114.35
670.0000000000,-114.30
671.0000000000,-114.25
672.0000000000,-114.20
673.0000000000,-114.16
674.0000000000,-114.14
675.0000000000,-114.12
676.0000000000,-114.08
677.0000000000,-114.03
678.0000000000,-113.99
679.0000000000,-113.94
680.0000000000,-113.89
681.0000000000,-113.85
682.0000000000,-113.80
683.0000000000,-113.75
684.0000000000,-113.70
685.0000000000,-113.66
686.0000000000,-113.61
687.0000000000,-113.56
688.0000000000,-113.51
689.0000000000,-113.47
690.0000000000,-113.42
691.0000000000,-113.37
692.0000000000,-113.33
693.0000000000,-113.28
694.0000000000,-113.24
695.0000000000,-113.19
696.0000000000,-113.14
697.0000000000,-113.10
698.0000000000,-113.05
699.0000000000,-113.01
700.0000000000,-112.96
701.0000000000,-112.91
702.0000000000,-112.87
703.0000000000,-112.82
704.0000000000,-112.78
705.0000000000,-112.73
706.0000000000,-112.68
707.0000000000,-112.64
708.0000000000,-112.59
709.0000000000,-112.55
710.0000000000,-112.50
711.0000000000,-112.46
712.0000000000,-112.41
713.0000000000,-112.37
714.0000000000,-112.32
715.0000000000,-112.27
716.0000000000,-112.23
717.0000000000,-112.18
718.0000000000,-112.14
719.0000000000,-112.10
720.0000000000,-112.05
721.0000000000,-112.01
722.0000000000,-111.96
723.0000000000,-111.92
724.0000000000,-111.87
725.0000000000,-111.83
726.0000000000,-111.78
727.0000000000,-111.75
728.0000000000,-111.71
729.0000000000,-111.67
730.0000000000,-111.62
731.0000000000,-111.58
732.0000000000,-111.54
733.0000000000,-111.50
734.0000000000,-111.46
735.0000000000,-111.42
736.0000000000,-111.37
737.0000000000,-111.33
738.0000000000,-111.29
739.0000000000,-111.24
740.0000000000,-111.21
741.0000000000,-111.16
742.0000000000,-111.12
743.0000000000,-111.08
744.0000000000,-111.03
745.0000000000,-110.99
746.0000000000,-110.95
747.0000000000,-110.90
748.0000000000,-110.86
749.0000000000,-110.82
750.0000000000,-110.78
751.0000000000,-110.73
752.0000000000,-110.69
753.0000000000,-110.66
754.0000000000,-110.61
755.0000000000,-110.57
756.0000000000,-110.53
757.0000000000,-110.49
758.0000000000,-110.44
759.0000000000,-110.40
760.0000000000,-110.36
761.0000000000,-110.32
762.0000000000,-110.28
763.0000000000,-110.24
764.0000000000,-110.20
765.0000000000,-110.16
766.0000000000,-110.12
767.0000000000,-110.08
768.0000000000,-110.03
769.0000000000,-109.99
770.0000000000,-109.95
771.0000000000,-109.91
772.0000000000,-109.87
773.0000000000,-109.82
774.0000000000,-109.78
775.0000000000,-109.74
776.0000000000,-109.70
777.0000000000,-109.66
778.0000000000,-109.62
779.0000000000,-109.58
780.0000000000,-109.53
781.0000000000,-109.49
782.0000000000,-109.45
783.0000000000,-109.41
784.0000000000,-109.37
785.0000000000,-109.33
786.0000000000,-109.29
787.0000000000,-109.25
788.0000000000,-109.20
789.0000000000,-109.17
790.0000000000,-109.13
791.0000000000,-109.08
792.0000000000,-109.04
793.0000000000,-109.00
794.0000000000,-108.97
795.0000000000,-108.93
796.0000000000,-108.89
797.0000000000,-108.85
798.0000000000,-108.81
799.0000000000,-108.77
800.0000000000,-108.73
801.0000000000,-108.69
802.0000000000,-108.65
803.0000000000,-108.61
804.0000000000,-108.57
805.0000000000,-108.53
806.0000000000,-108.49
807.0000000000,-108.45
808.0000000000,-108.41
809.0000000000,-108.38
810.0000000000,-108.36
811.0000000000,-108.34
812.0000000000,-108.31
813.0000000000,-108.27
814.0000000000,-108.23
815.0000000000,-108.19
816.0000000000,-108.15
817.0000000000,-108.12
818.0000000000,-108.08
819.0000000000,-108.04
820.0000000000,-108.00
821.0000000000,-107.96
822.0000000000,-107.92
823.0000000000,-107.88
824.0000000000,-107.84
825.0000000000,-107.80
826.0000000000,-107.76
827.0000000000,-107.73
828.0000000000,-107.69
829.0000000000,-107.65
830.0000000000,-107.61
831.0000000000,-107.57
832.0000000000,-107.54
833.0000000000,-107.51
834.0000000000,-107.47
835.0000000000,-107.44
836.0000000000,-107.40
837.0000000000,-107.37
838.0000000000,-107.34
839.0000000000,-107.30
840.0000000000,-107.26
841.0000000000,-107.23
842.0000000000,-107.19
843.0000000000,-107.15
844.0000000000,-107.12
845.0000000000,-107.08
846.0000000000,-107.04
847.0000000000,-107.01
848.0000000000,-106.98
849.0000000000,-106.94
850.0000000000,-106.90
851.0000000000,-106.87
852.0000000000,-106.83
853.0000000000,-106.79
854.0000000000,-106.75
855.0000000000,-106.72
856.0000000000,-106.68
857.0000000000,-106.64
858.0000000000,-106.60
859.0000000000,-106.57
860.0000000000,-106.53
861.0000000000,-106.52
862.0000000000,-106.51
863.0000000000,-106.50
864.0000000000,-106.47
865.0000000000,-106.44
866.0000000000,-106.42
867.0000000000,-106.41
868.0000000000,-106.38
869.0000000000,-106.34
870.0000000000,-106.31
871.0000000000,-106.28
872.0000000000,-106.25
873.0000000000,-106.21
874.0000000000,-106.18
875.0000000000,-106.15
876.0000000000,-106.11
877.0000000000,-106.08
878.0000000000,-106.04
879.0000000000,-106.03
880.0000000000,-106.00
881.0000000000,-105.98
882.0000000000,-105.95
883.0000000000,-105.92
884.0000000000,-105.88
885.0000000000,-105.85
886.0000000000,-105.81
887.0000000000,-105.77
888.0000000000,-105.74
889.0000000000,-105.70
890.0000000000,-105.67
891.0000000000,-105.63
892.0000000000,-105.59
893.0000000000,-105.56
894.0000000000,-105.52
895.0000000000,-105.50
896.0000000000,-105.47
897.0000000000,-105.45
898.0000000000,-105.42
899.0000000000,-105.38
900.0000000000,-105.35
901.0000000000,-105.32
902.0000000000,-105.29
903.0000000000,-105.25
904.0000000000,-105.22
905.0000000000,-105.19
906.0000000000,-105.15
907.0000000000,-105.12
908.0000000000,-105.09
909.0000000000,-105.07
910.0000000000,-105.03
911.0000000000,-105.00
912.0000000000,-104.97
913.0000000000,-104.93
914.0000000000,-104.90
915.0000000000,-104.86
916.0000000000,-104.83
917.0000000000,-104.79
918.0000000000,-104.76
919.0000000000,-104.73
920.0000000000,-104.70
921.0000000000,-104.67
922.0000000000,-104.63
923.0000000000,-104.60
924.0000000000,-104.56
925.0000000000,-104.53
926.0000000000,-104.49
927.0000000000,-104.46
928.0000000000,-104.43
929.0000000000,-104.39
930.0000000000,-104.36
931.0000000000,-104.32
932.0000000000,-104.29
933.0000000000,-104.25
934.0000000000,-104.22
935.0000000000,-104.19
936.0000000000,-104.15
937.0000000000,-104.12
938.0000000000,-104.08
939.0000000000,-104.05
940.0000000000,-104.02
941.0000000000,-103.98
942.0000000000,-103.95
943.0000000000,-103.92
944.0000000000,-103.89
945.0000000000,-103.85
946.0000000000,-103.82
947.0000000000,-103.79
948.0000000000,-103.75
949.0000000000,-103.72
950.0000000000,-103.69
951.0000000000,-103.65
952.0000000000,-103.62
953.0000000000,-103.59
954.0000000000,-103.55
955.0000000000,-103.52
956.0000000000,-103.49
957.0000000000,-103.46
958.0000000000,-103.44
959.0000000000,-103.41
960.0000000000,-103.38
961.0000000000,-103.34
962.0000000000,-103.32
963.0000000000,-103.29
964.0000000000,-103.26
965.0000000000,-103.23
966.0000000000,-103.19
967.0000000000,-103.16
968.0000000000,-103.13
969.0000000000,-103.10
970.0000000000,-103.07
971.0000000000,-103.04
972.0000000000,-103.00
973.0000000000,-102.97
974.0000000000,-102.94
975.0000000000,-102.91
976.0000000000,-102.88
977.0000000000,-102.84
978.0000000000,-102.81
979.0000000000,-102.78
980.0000000000,-102.75
981.0000000000,-102.71
982.0000000000,-102.68
983.0000000000,-102.66
984.0000000000,-102.62
985.0000000000,-102.60
986.0000000000,-102.56
987.0000000000,-102.53
988.0000000000,-102.50
989.0000000000,-102.47
990.0000000000,-102.44
991.0000000000,-102.41
992.0000000000,-102.37
993.0000000000,-102.34
994.0000000000,-102.31
995.0000000000,-102.28
996.0000000000,-102.25
997.0000000000,-102.22
998.0000000000,-102.19
999.0000000000,-102.15
1000.000000000,-102.12
1001.000000000,-102.09
1002.000000000,-102.06
1003.000000000,-102.03
1004.000000000,-102.00
1005.000000000,-101.97
1006.000000000,-101.94
1007.000000000,-101.91
1008.000000000,-101.88
1009.000000000,-101.85
1010.000000000,-101.81
1011.000000000,-101.78
1012.000000000,-101.77
1013.000000000,-101.75
1014.000000000,-101.72
1015.000000000,-101.69
1016.000000000,-101.66
1017.000000000,-101.63
1018.000000000,-101.60
1019.000000000,-101.57
1020.000000000,-101.54
1021.000000000,-101.51
1022.000000000,-101.48
1023.000000000,-101.45
1024.000000000,-101.42
1025.000000000,-101.39
1026.000000000,-101.36
1027.000000000,-101.38
1028.000000000,-101.38
1029.000000000,-101.36
1030.000000000,-101.33
1031.000000000,-101.30
1032.000000000,-101.27
1033.000000000,-101.25
1034.000000000,-101.24
1035.000000000,-101.22
1036.000000000,-101.19
1037.000000000,-101.16
1038.000000000,-101.13
1039.000000000,-101.10
1040.000000000,-101.07
1041.000000000,-101.04
1042.000000000,-101.01
1043.000000000,-100.99
1044.000000000,-100.96
1045.000000000,-100.93
1046.000000000,-100.90
1047.000000000,-100.87
1048.000000000,-100.84
1049.000000000,-100.81
1050.000000000,-100.78
1051.000000000,-100.75
1052.000000000,-100.72
1053.000000000,-100.69
1054.000000000,-100.67
1055.000000000,-100.64
1056.000000000,-100.61
1057.000000000,-100.58
1058.000000000,-100.55
1059.000000000,-100.52
1060.000000000,-100.49
1061.000000000,-100.47
1062.000000000,-100.45
1063.000000000,-100.43
1064.000000000,-100.40
1065.000000000,-100.37
1066.000000000,-100.35
1067.000000000,-100.32
1068.000000000,-100.29
1069.000000000,-100.26
1070.000000000,-100.23
1071.000000000,-100.20
1072.000000000,-100.17
1073.000000000,-100.14
1074.000000000,-100.12
1075.000000000,-100.09
1076.000000000,-100.06
1077.000000000,-100.05
1078.000000000,-100.02
1079.000000000,-99.997
1080.000000000,-99.970
1081.000000000,-99.942
1082.000000000,-99.913
1083.000000000,-99.885
1084.000000000,-99.857
1085.000000000,-99.828
1086.000000000,-99.800
1087.000000000,-99.772
1088.000000000,-99.744
1089.000000000,-99.715
1090.000000000,-99.687
1091.000000000,-99.675
1092.000000000,-99.654
1093.000000000,-99.628
1094.000000000,-99.601
1095.000000000,-99.574
1096.000000000,-99.546
1097.000000000,-99.519
1098.000000000,-99.494
1099.000000000,-99.467
1100.000000000,-99.439
1101.000000000,-99.411
1102.000000000,-99.384
1103.000000000,-99.356
1104.000000000,-99.328
1105.000000000,-99.301
1106.000000000,-99.273
1107.000000000,-99.246
1108.000000000,-99.218
1109.000000000,-99.191
1110.000000000,-99.163
1111.000000000,-99.136
1112.000000000,-99.108
1113.000000000,-99.081
1114.000000000,-99.054
1115.000000000,-99.026
1116.000000000,-98.999
1117.000000000,-98.972
1118.000000000,-98.945
1119.000000000,-98.918
1120.000000000,-98.891
1121.000000000,-98.864
1122.000000000,-98.846
1123.000000000,-98.822
1124.000000000,-98.796
1125.000000000,-98.769
1126.000000000,-98.743
1127.000000000,-98.716
1128.000000000,-98.689
1129.000000000,-98.662
1130.000000000,-98.635
1131.000000000,-98.609
1132.000000000,-98.582
1133.000000000,-98.555
1134.000000000,-98.529
1135.000000000,-98.502
1136.000000000,-98.476
1137.000000000,-98.449
1138.000000000,-98.423
1139.000000000,-98.396
1140.000000000,-98.370
1141.000000000,-98.344
1142.000000000,-98.317
1143.000000000,-98.291
1144.000000000,-98.265
1145.000000000,-98.239
1146.000000000,-98.212
1147.000000000,-98.186
1148.000000000,-98.164
1149.000000000,-98.149
1150.000000000,-98.126
1151.000000000,-98.101
1152.000000000,-98.075
1153.000000000,-98.049
1154.000000000,-98.024
1155.000000000,-97.998
1156.000000000,-97.972
1157.000000000,-97.946
1158.000000000,-97.920
1159.000000000,-97.894
1160.000000000,-97.869
1161.000000000,-97.843
1162.000000000,-97.817
1163.000000000,-97.809
1164.000000000,-97.798
1165.000000000,-97.793
1166.000000000,-97.789
1167.000000000,-97.779
1168.000000000,-97.759
1169.000000000,-97.735
1170.000000000,-97.710
1171.000000000,-97.685
1172.000000000,-97.660
1173.000000000,-97.635
1174.000000000,-97.617
1175.000000000,-97.594
1176.000000000,-97.569
1177.000000000,-97.544
1178.000000000,-97.519
1179.000000000,-97.494
1180.000000000,-97.469
1181.000000000,-97.444
1182.000000000,-97.419
1183.000000000,-97.394
1184.000000000,-97.369
1185.000000000,-97.344
1186.000000000,-97.319
1187.000000000,-97.294
1188.000000000,-97.269
1189.000000000,-97.244
1190.000000000,-97.219
1191.000000000,-97.194
1192.000000000,-97.169
1193.000000000,-97.144
1194.000000000,-97.119
1195.000000000,-97.095
1196.000000000,-97.070
1197.000000000,-97.045
1198.000000000,-97.021
1199.000000000,-97.003
1200.000000000,-96.980
1201.000000000,-96.956
1202.000000000,-96.932
1203.000000000,-96.955
1204.000000000,-96.951
1205.000000000,-96.934
1206.000000000,-96.913
1207.000000000,-96.890
1208.000000000,-96.866
1209.000000000,-96.842
1210.000000000,-96.818
1211.000000000,-96.794
1212.000000000,-96.770
1213.000000000,-96.750
1214.000000000,-96.727
1215.000000000,-96.703
1216.000000000,-96.679
1217.000000000,-96.655
1218.000000000,-96.631
1219.000000000,-96.607
1220.000000000,-96.582
1221.000000000,-96.558
1222.000000000,-96.534
1223.000000000,-96.510
1224.000000000,-96.486
1225.000000000,-96.464
1226.000000000,-96.440
1227.000000000,-96.416
1228.000000000,-96.392
1229.000000000,-96.369
1230.000000000,-96.345
1231.000000000,-96.324
1232.000000000,-96.302
1233.000000000,-96.279
1234.000000000,-96.261
1235.000000000,-96.254
1236.000000000,-96.237
1237.000000000,-96.216
1238.000000000,-96.193
1239.000000000,-96.170
1240.000000000,-96.147
1241.000000000,-96.123
1242.000000000,-96.100
1243.000000000,-96.076
1244.000000000,-96.053
1245.000000000,-96.029
1246.000000000,-96.007
1247.000000000,-95.983
1248.000000000,-95.962
1249.000000000,-95.969
1250.000000000,-95.960
1251.000000000,-95.942
1252.000000000,-95.921
1253.000000000,-95.898
1254.000000000,-95.876
1255.000000000,-95.852
1256.000000000,-95.829
1257.000000000,-95.806
1258.000000000,-95.783
1259.000000000,-95.760
1260.000000000,-95.737
1261.000000000,-95.714
1262.000000000,-95.691
1263.000000000,-95.668
1264.000000000,-95.645
1265.000000000,-95.622
1266.000000000,-95.599
1267.000000000,-95.583
1268.000000000,-95.562
1269.000000000,-95.540
1270.000000000,-95.517
1271.000000000,-95.495
1272.000000000,-95.472
1273.000000000,-95.456
1274.000000000,-95.485
1275.000000000,-95.477
1276.000000000,-95.460
1277.000000000,-95.440
1278.000000000,-95.419
1279.000000000,-95.397
1280.000000000,-95.374
1281.000000000,-95.352
1282.000000000,-95.329
1283.000000000,-95.306
1284.000000000,-95.284
1285.000000000,-95.261
1286.000000000,-95.239
1287.000000000,-95.216
1288.000000000,-95.194
1289.000000000,-95.172
1290.000000000,-95.149
1291.000000000,-95.127
1292.000000000,-95.105
1293.000000000,-95.082
1294.000000000,-95.060
1295.000000000,-95.038
1296.000000000,-95.016
1297.000000000,-94.994
1298.000000000,-94.971
1299.000000000,-94.949
1300.000000000,-94.927
1301.000000000,-94.905
1302.000000000,-94.883
1303.000000000,-94.861
1304.000000000,-94.845
1305.000000000,-94.825
1306.000000000,-94.803
1307.000000000,-94.782
1308.000000000,-94.760
1309.000000000,-94.739
1310.000000000,-94.717
1311.000000000,-94.695
1312.000000000,-94.674
1313.000000000,-94.652
1314.000000000,-94.630
1315.000000000,-94.609
1316.000000000,-94.587
1317.000000000,-94.565
1318.000000000,-94.544
1319.000000000,-94.522
1320.000000000,-94.501
1321.000000000,-94.498
1322.000000000,-94.497
1323.000000000,-94.487
1324.000000000,-94.471
1325.000000000,-94.462
1326.000000000,-94.448
1327.000000000,-94.430
1328.000000000,-94.449
1329.000000000,-94.442
1330.000000000,-94.433
1331.000000000,-94.425
1332.000000000,-94.408
1333.000000000,-94.389
1334.000000000,-94.369
1335.000000000,-94.348
1336.000000000,-94.328
1337.000000000,-94.309
1338.000000000,-94.290
1339.000000000,-94.272
1340.000000000,-94.254
1341.000000000,-94.235
1342.000000000,-94.220
1343.000000000,-94.201
1344.000000000,-94.180
1345.000000000,-94.160
1346.000000000,-94.139
1347.000000000,-94.118
1348.000000000,-94.097
1349.000000000,-94.076
1350.000000000,-94.057
1351.000000000,-94.037
1352.000000000,-94.021
1353.000000000,-94.002
1354.000000000,-93.984
1355.000000000,-93.964
1356.000000000,-93.943
1357.000000000,-93.923
1358.000000000,-93.902
1359.000000000,-93.881
1360.000000000,-93.861
1361.000000000,-93.840
1362.000000000,-93.819
1363.000000000,-93.799
1364.000000000,-93.803
1365.000000000,-93.844
1366.000000000,-93.845
1367.000000000,-93.832
1368.000000000,-93.815
1369.000000000,-93.796
1370.000000000,-93.776
1371.000000000,-93.756
1372.000000000,-93.735
1373.000000000,-93.715
1374.000000000,-93.694
1375.000000000,-93.674
1376.000000000,-93.654
1377.000000000,-93.633
1378.000000000,-93.613
1379.000000000,-93.593
1380.000000000,-93.572
1381.000000000,-93.552
1382.000000000,-93.532
1383.000000000,-93.511
1384.000000000,-93.491
1385.000000000,-93.471
1386.000000000,-93.451
1387.000000000,-93.431
1388.000000000,-93.410
1389.000000000,-93.390
1390.000000000,-93.370
1391.000000000,-93.350
1392.000000000,-93.330
1393.000000000,-93.310
1394.000000000,-93.290
1395.000000000,-93.270
1396.000000000,-93.251
1397.000000000,-93.231
1398.000000000,-93.211
1399.000000000,-93.191
1400.000000000,-93.171
1401.000000000,-93.151
1402.000000000,-93.131
1403.000000000,-93.112
1404.000000000,-93.103
1405.000000000,-93.086
1406.000000000,-93.067
1407.000000000,-93.050
1408.000000000,-93.031
1409.000000000,-93.011
1410.000000000,-93.008
1411.000000000,-92.992
1412.000000000,-92.975
1413.000000000,-92.956
1414.000000000,-92.937
1415.000000000,-92.917
1416.000000000,-92.898
1417.000000000,-92.878
1418.000000000,-92.859
1419.000000000,-92.839
1420.000000000,-92.820
1421.000000000,-92.801
1422.000000000,-92.781
1423.000000000,-92.762
1424.000000000,-92.743
1425.000000000,-92.723
1426.000000000,-92.705
1427.000000000,-92.687
1428.000000000,-92.667
1429.000000000,-92.648
1430.000000000,-92.629
1431.000000000,-92.610
1432.000000000,-92.591
1433.000000000,-92.578
1434.000000000,-92.571
1435.000000000,-92.590
1436.000000000,-92.583
1437.000000000,-92.569
1438.000000000,-92.552
1439.000000000,-92.534
1440.000000000,-92.515
1441.000000000,-92.496
1442.000000000,-92.477
1443.000000000,-92.459
1444.000000000,-92.441
1445.000000000,-92.422
1446.000000000,-92.403
1447.000000000,-92.384
1448.000000000,-92.365
1449.000000000,-92.346
1450.000000000,-92.327
1451.000000000,-92.309
1452.000000000,-92.291
1453.000000000,-92.272
1454.000000000,-92.255
1455.000000000,-92.237
1456.000000000,-92.218
1457.000000000,-92.199
1458.000000000,-92.181
1459.000000000,-92.162
1460.000000000,-92.144
1461.000000000,-92.126
1462.000000000,-92.107
1463.000000000,-92.089
1464.000000000,-92.071
1465.000000000,-92.053
1466.000000000,-92.034
1467.000000000,-92.016
1468.000000000,-91.998
1469.000000000,-91.979
1470.000000000,-91.961
1471.000000000,-91.943
1472.000000000,-91.924
1473.000000000,-91.906
1474.000000000,-91.888
1475.000000000,-91.871
1476.000000000,-91.856
1477.000000000,-91.844
1478.000000000,-91.827
1479.000000000,-91.817
1480.000000000,-91.801
1481.000000000,-91.784
1482.000000000,-91.766
1483.000000000,-91.748
1484.000000000,-91.730
1485.000000000,-91.712
1486.000000000,-91.694
1487.000000000,-91.676
1488.000000000,-91.658
1489.000000000,-91.641
1490.000000000,-91.623
1491.000000000,-91.605
1492.000000000,-91.587
1493.000000000,-91.569
1494.000000000,-91.552
1495.000000000,-91.534
1496.000000000,-91.516
1497.000000000,-91.498
1498.000000000,-91.481
1499.000000000,-91.463
1500.000000000,-91.445
1501.000000000,-91.428
1502.000000000,-91.410
1503.000000000,-91.392
1504.000000000,-91.375
1505.000000000,-91.357
1506.000000000,-91.363
1507.000000000,-91.351
1508.000000000,-91.336
1509.000000000,-91.320
1510.000000000,-91.303
1511.000000000,-91.286
1512.000000000,-91.271
1513.000000000,-91.255
1514.000000000,-91.237
1515.000000000,-91.220
1516.000000000,-91.203
1517.000000000,-91.185
1518.000000000,-91.168
1519.000000000,-91.151
1520.000000000,-91.133
1521.000000000,-91.116
1522.000000000,-91.099
1523.000000000,-91.081
1524.000000000,-91.064
1525.000000000,-91.049
1526.000000000,-91.032
1527.000000000,-91.015
1528.000000000,-90.998
1529.000000000,-90.981
1530.000000000,-90.963
1531.000000000,-90.947
1532.000000000,-90.930
1533.000000000,-90.913
1534.000000000,-90.896
1535.000000000,-90.879
1536.000000000,-90.862
1537.000000000,-90.845
1538.000000000,-90.828
1539.000000000,-90.811
1540.000000000,-90.794
1541.000000000,-90.777
1542.000000000,-90.760
1543.000000000,-90.744
1544.000000000,-90.727
1545.000000000,-90.710
1546.000000000,-90.694
1547.000000000,-90.677
1548.000000000,-90.660
1549.000000000,-90.654
1550.000000000,-90.640
1551.000000000,-90.624
1552.000000000,-90.608
1553.000000000,-90.611
1554.000000000,-90.599
1555.000000000,-90.584
1556.000000000,-90.569
1557.000000000,-90.553
1558.000000000,-90.536
1559.000000000,-90.520
1560.000000000,-90.503
1561.000000000,-90.486
1562.000000000,-90.476
1563.000000000,-90.463
1564.000000000,-90.450
1565.000000000,-90.443
1566.000000000,-90.429
1567.000000000,-90.414
1568.000000000,-90.401
1569.000000000,-90.386
1570.000000000,-90.370
1571.000000000,-90.354
1572.000000000,-90.337
1573.000000000,-90.321
1574.000000000,-90.305
1575.000000000,-90.288
1576.000000000,-90.272
1577.000000000,-90.256
1578.000000000,-90.240
1579.000000000,-90.223
1580.000000000,-90.207
1581.000000000,-90.191
1582.000000000,-90.175
1583.000000000,-90.159
1584.000000000,-90.143
1585.000000000,-90.126
1586.000000000,-90.110
1587.000000000,-90.094
1588.000000000,-90.078
1589.000000000,-90.062
1590.000000000,-90.046
1591.000000000,-90.030
1592.000000000,-90.022
1593.000000000,-90.008
1594.000000000,-89.993
1595.000000000,-89.978
1596.000000000,-89.962
1597.000000000,-89.946
1598.000000000,-89.931
1599.000000000,-89.915
1600.000000000,-89.899
1601.000000000,-89.899
1602.000000000,-89.888
1603.000000000,-89.887
1604.000000000,-89.876
1605.000000000,-89.862
1606.000000000,-89.847
1607.000000000,-89.832
1608.000000000,-89.816
1609.000000000,-89.801
1610.000000000,-89.801
1611.000000000,-89.789
1612.000000000,-89.828
1613.000000000,-89.831
1614.000000000,-89.824
1615.000000000,-89.815
1616.000000000,-89.811
1617.000000000,-89.799
1618.000000000,-89.785
1619.000000000,-89.770
1620.000000000,-89.755
1621.000000000,-89.739
1622.000000000,-89.723
1623.000000000,-89.707
1624.000000000,-89.692
1625.000000000,-89.676
1626.000000000,-89.660
1627.000000000,-89.645
1628.000000000,-89.629
1629.000000000,-89.614
1630.000000000,-89.598
1631.000000000,-89.583
1632.000000000,-89.567
1633.000000000,-89.552
1634.000000000,-89.536
1635.000000000,-89.521
1636.000000000,-89.506
1637.000000000,-89.490
1638.000000000,-89.475
1639.000000000,-89.464
1640.000000000,-89.451
1641.000000000,-89.436
1642.000000000,-89.421
1643.000000000,-89.406
1644.000000000,-89.391
1645.000000000,-89.376
1646.000000000,-89.360
1647.000000000,-89.346
1648.000000000,-89.331
1649.000000000,-89.322
1650.000000000,-89.317
1651.000000000,-89.304
1652.000000000,-89.290
1653.000000000,-89.275
1654.000000000,-89.260
1655.000000000,-89.245
1656.000000000,-89.232
1657.000000000,-89.220
1658.000000000,-89.210
1659.000000000,-89.198
1660.000000000,-89.185
1661.000000000,-89.172
1662.000000000,-89.157
1663.000000000,-89.142
1664.000000000,-89.128
1665.000000000,-89.113
1666.000000000,-89.113
1667.000000000,-89.102
1668.000000000,-89.089
1669.000000000,-89.074
1670.000000000,-89.060
1671.000000000,-89.045
1672.000000000,-89.030
1673.000000000,-89.017
1674.000000000,-89.004
1675.000000000,-88.992
1676.000000000,-88.981
1677.000000000,-88.967
1678.000000000,-88.953
1679.000000000,-88.939
1680.000000000,-88.924
1681.000000000,-88.911
1682.000000000,-88.916
1683.000000000,-88.906
1684.000000000,-88.894
1685.000000000,-88.880
1686.000000000,-88.866
1687.000000000,-88.851
1688.000000000,-88.837
1689.000000000,-88.823
1690.000000000,-88.810
1691.000000000,-88.796
1692.000000000,-88.781
1693.000000000,-88.767
1694.000000000,-88.752
1695.000000000,-88.738
1696.000000000,-88.723
1697.000000000,-88.714
1698.000000000,-88.706
1699.000000000,-88.694
1700.000000000,-88.685
1701.000000000,-88.672
1702.000000000,-88.658
1703.000000000,-88.644
1704.000000000,-88.629
1705.000000000,-88.615
1706.000000000,-88.601
1707.000000000,-88.587
1708.000000000,-88.572
1709.000000000,-88.558
1710.000000000,-88.544
1711.000000000,-88.530
1712.000000000,-88.516
1713.000000000,-88.501
1714.000000000,-88.487
1715.000000000,-88.473
1716.000000000,-88.459
1717.000000000,-88.445
1718.000000000,-88.431
1719.000000000,-88.417
1720.000000000,-88.403
1721.000000000,-88.388
1722.000000000,-88.374
1723.000000000,-88.360
1724.000000000,-88.347
1725.000000000,-88.333
1726.000000000,-88.319
1727.000000000,-88.305
1728.000000000,-88.291
1729.000000000,-88.295
1730.000000000,-88.295
1731.000000000,-88.319
1732.000000000,-88.349
1733.000000000,-88.363
1734.000000000,-88.363
1735.000000000,-88.355
1736.000000000,-88.344
1737.000000000,-88.331
1738.000000000,-88.327
1739.000000000,-88.317
1740.000000000,-88.305
1741.000000000,-88.291
1742.000000000,-88.278
1743.000000000,-88.264
1744.000000000,-88.255
1745.000000000,-88.243
1746.000000000,-88.229
1747.000000000,-88.216
1748.000000000,-88.202
1749.000000000,-88.188
1750.000000000,-88.175
1751.000000000,-88.161
1752.000000000,-88.147
1753.000000000,-88.133
1754.000000000,-88.120
1755.000000000,-88.106
1756.000000000,-88.092
1757.000000000,-88.078
1758.000000000,-88.065
1759.000000000,-88.051
1760.000000000,-88.038
1761.000000000,-88.024
1762.000000000,-88.010
1763.000000000,-87.997
1764.000000000,-87.983
1765.000000000,-87.970
1766.000000000,-87.956
1767.000000000,-87.943
1768.000000000,-87.929
1769.000000000,-87.916
1770.000000000,-87.902
1771.000000000,-87.889
1772.000000000,-87.875
1773.000000000,-87.862
1774.000000000,-87.848
1775.000000000,-87.835
1776.000000000,-87.822
1777.000000000,-87.810
1778.000000000,-87.797
1779.000000000,-87.784
1780.000000000,-87.771
1781.000000000,-87.758
1782.000000000,-87.745
1783.000000000,-87.731
1784.000000000,-87.718
1785.000000000,-87.705
1786.000000000,-87.691
1787.000000000,-87.678
1788.000000000,-87.665
1789.000000000,-87.652
1790.000000000,-87.639
1791.000000000,-87.626
1792.000000000,-87.612
1793.000000000,-87.599
1794.000000000,-87.586
1795.000000000,-87.573
1796.000000000,-87.560
1797.000000000,-87.547
1798.000000000,-87.534
1799.000000000,-87.521
1800.000000000,-87.508
1801.000000000,-87.499
1802.000000000,-87.504
1803.000000000,-87.500
1804.000000000,-87.490
1805.000000000,-87.478
1806.000000000,-87.466
1807.000000000,-87.453
1808.000000000,-87.440
1809.000000000,-87.427
1810.000000000,-87.414
1811.000000000,-87.402
1812.000000000,-87.395
1813.000000000,-87.384
1814.000000000,-87.373
1815.000000000,-87.361
1816.000000000,-87.348
1817.000000000,-87.335
1818.000000000,-87.322
1819.000000000,-87.310
1820.000000000,-87.297
1821.000000000,-87.284
1822.000000000,-87.272
1823.000000000,-87.260
1824.000000000,-87.247
1825.000000000,-87.235
1826.000000000,-87.222
1827.000000000,-87.209
1828.000000000,-87.197
1829.000000000,-87.184
1830.000000000,-87.171
1831.000000000,-87.159
1832.000000000,-87.146
1833.000000000,-87.133
1834.000000000,-87.121
1835.000000000,-87.108
1836.000000000,-87.096
1837.000000000,-87.083
1838.000000000,-87.071
1839.000000000,-87.058
1840.000000000,-87.046
1841.000000000,-87.033
1842.000000000,-87.021
1843.000000000,-87.009
1844.000000000,-86.996
1845.000000000,-86.984
1846.000000000,-86.972
1847.000000000,-86.959
1848.000000000,-86.947
1849.000000000,-86.935
1850.000000000,-86.922
1851.000000000,-86.910
1852.000000000,-86.898
1853.000000000,-86.885
1854.000000000,-86.873
1855.000000000,-86.861
1856.000000000,-86.849
1857.000000000,-86.836
1858.000000000,-86.824
1859.000000000,-86.812
1860.000000000,-86.800
1861.000000000,-86.788
1862.000000000,-86.776
1863.000000000,-86.764
1864.000000000,-86.752
1865.000000000,-86.739
1866.000000000,-86.727
1867.000000000,-86.715
1868.000000000,-86.703
1869.000000000,-86.691
1870.000000000,-86.680
1871.000000000,-86.669
1872.000000000,-86.657
1873.000000000,-86.645
1874.000000000,-86.633
1875.000000000,-86.621
1876.000000000,-86.611
1877.000000000,-86.604
1878.000000000,-86.613
1879.000000000,-86.607
1880.000000000,-86.598
1881.000000000,-86.587
1882.000000000,-86.576
1883.000000000,-86.564
1884.000000000,-86.552
1885.000000000,-86.541
1886.000000000,-86.530
1887.000000000,-86.518
1888.000000000,-86.506
1889.000000000,-86.494
1890.000000000,-86.482
1891.000000000,-86.471
1892.000000000,-86.459
1893.000000000,-86.447
1894.000000000,-86.435
1895.000000000,-86.423
1896.000000000,-86.411
1897.000000000,-86.400
1898.000000000,-86.388
1899.000000000,-86.376
1900.000000000,-86.364
1901.000000000,-86.353
1902.000000000,-86.341
1903.000000000,-86.329
1904.000000000,-86.318
1905.000000000,-86.306
1906.000000000,-86.294
1907.000000000,-86.283
1908.000000000,-86.271
1909.000000000,-86.260
1910.000000000,-86.248
1911.000000000,-86.236
1912.000000000,-86.225
1913.000000000,-86.214
1914.000000000,-86.203
1915.000000000,-86.192
1916.000000000,-86.180
1917.000000000,-86.169
1918.000000000,-86.157
1919.000000000,-86.146
1920.000000000,-86.134
1921.000000000,-86.123
1922.000000000,-86.111
1923.000000000,-86.100
1924.000000000,-86.089
1925.000000000,-86.077
1926.000000000,-86.066
1927.000000000,-86.055
1928.000000000,-86.043
1929.000000000,-86.032
1930.000000000,-86.021
1931.000000000,-86.010
1932.000000000,-85.999
1933.000000000,-85.987
1934.000000000,-85.976
1935.000000000,-85.965
1936.000000000,-85.954
1937.000000000,-85.943
1938.000000000,-85.932
1939.000000000,-85.921
1940.000000000,-85.909
1941.000000000,-85.898
1942.000000000,-85.890
1943.000000000,-85.880
1944.000000000,-85.869
1945.000000000,-85.858
1946.000000000,-85.847
1947.000000000,-85.836
1948.000000000,-85.825
1949.000000000,-85.815
1950.000000000,-85.826
1951.000000000,-85.824
1952.000000000,-85.816
1953.000000000,-85.806
1954.000000000,-85.796
1955.000000000,-85.785
1956.000000000,-85.774
1957.000000000,-85.763
1958.000000000,-85.752
1959.000000000,-85.741
1960.000000000,-85.730
1961.000000000,-85.719
1962.000000000,-85.708
1963.000000000,-85.697
1964.000000000,-85.686
1965.000000000,-85.675
1966.000000000,-85.666
1967.000000000,-85.677
1968.000000000,-85.672
1969.000000000,-85.663
1970.000000000,-85.653
1971.000000000,-85.643
1972.000000000,-85.632
1973.000000000,-85.621
1974.000000000,-85.610
1975.000000000,-85.600
1976.000000000,-85.589
1977.000000000,-85.578
1978.000000000,-85.567
1979.000000000,-85.556
1980.000000000,-85.545
1981.000000000,-85.536
1982.000000000,-85.525
1983.000000000,-85.515
1984.000000000,-85.504
1985.000000000,-85.493
1986.000000000,-85.482
1987.000000000,-85.472
1988.000000000,-85.461
1989.000000000,-85.450
1990.000000000,-85.440
1991.000000000,-85.429
1992.000000000,-85.418
1993.000000000,-85.408
1994.000000000,-85.397
1995.000000000,-85.387
1996.000000000,-85.378
1997.000000000,-85.367
1998.000000000,-85.357
1999.000000000,-85.347
2000.000000000,-85.336
2001.000000000,-85.326
2002.000000000,-85.315
2003.000000000,-85.305
2004.000000000,-85.294
2005.000000000,-85.284
2006.000000000,-85.273
2007.000000000,-85.264
2008.000000000,-85.254
2009.000000000,-85.244
2010.000000000,-85.233
2011.000000000,-85.223
2012.000000000,-85.215
2013.000000000,-85.209
2014.000000000,-85.208
2015.000000000,-85.210
2016.000000000,-85.207
2017.000000000,-85.206
2018.000000000,-85.198
2019.000000000,-85.189
2020.000000000,-85.179
2021.000000000,-85.169
2022.000000000,-85.159
2023.000000000,-85.148
2024.000000000,-85.138
2025.000000000,-85.128
2026.000000000,-85.117
2027.000000000,-85.107
2028.000000000,-85.097
2029.000000000,-85.086
2030.000000000,-85.076
2031.000000000,-85.066
2032.000000000,-85.056
2033.000000000,-85.045
2034.000000000,-85.035
2035.000000000,-85.025
2036.000000000,-85.015
2037.000000000,-85.005
2038.000000000,-85.016
2039.000000000,-85.011
2040.000000000,-85.004
2041.000000000,-84.995
2042.000000000,-84.985
2043.000000000,-84.975
2044.000000000,-84.965
2045.000000000,-84.955
2046.000000000,-84.945
2047.000000000,-84.935
2048.000000000,-84.925
2049.000000000,-84.923
2050.000000000,-84.920
2051.000000000,-84.920
2052.000000000,-84.914
2053.000000000,-84.906
2054.000000000,-84.897
2055.000000000,-84.887
2056.000000000,-84.877
2057.000000000,-84.867
2058.000000000,-84.859
2059.000000000,-84.852
2060.000000000,-84.843
2061.000000000,-84.834
2062.000000000,-84.824
2063.000000000,-84.814
2064.000000000,-84.804
2065.000000000,-84.794
2066.000000000,-84.784
2067.000000000,-84.774
2068.000000000,-84.764
2069.000000000,-84.754
