time,RECHARGE,RECHARGE,RECHARGE,RECHARGE,RECHARGE,RECHARGE,RECHARGE,RECHARGE,RECHARGE,RECHARGE,RECHARGE,RECHARGE,DISCHARGE,DISCHARGE,DISCHARGE,DISCHARGE,DISCHARGE,DISCHARGE,DISCHARGE,DISCHARGE,DISCHARGE,DISCHARGE,DISCHARGE,DISCHARGE,INFILT,INFILT,INFILT,INFILT,INFILT,INFILT,INFILT,INFILT,INFILT,INFILT,INFILT,INFILT,REJINFILT,REJINFILT,REJINFILT,REJINFILT,REJINFILT,REJINFILT,REJINFILT,REJINFILT,REJINFILT,REJINFILT,REJINFILT,REJINFILT
1.000000000000,0.62679E+07,0.12107E+07,0.20314E+07,0.18706E+07,0.19212E+07,0.16609E+07,0.29613E+07,0.31281E+06,0.23273E+07,0.39805E+06,0.11042E+07,0.65871E+06,0.0000,-19173.,-13409.,-3024.4,-4746.3,-10089.,-32014.,-992.56,-34832.,-11175.,-13574.,-2771.4,61.694,169.16,159.41,95.785,70.442,127.51,115.89,53.083,253.98,104.81,165.29,96.039,0.0000,-20.300,-9.2034,-2.9731,-2.5888,-2.7198,-16.664,-2.4438,-26.525,-19.721,-10.791,-22.621
2.000000000000,0.59483E+07,0.75995E+06,0.10705E+07,0.11206E+07,0.13102E+07,0.63229E+06,0.18395E+07,0.25182E+06,0.94509E+06,0.15684E+06,0.38829E+06,0.38977E+06,0.0000,-20932.,-12946.,-3006.2,-4639.0,-9846.9,-33390.,-832.48,-34649.,-11143.,-15045.,-2294.9,7.6246,271.62,247.67,101.11,36.729,185.13,194.85,0.0000,662.94,177.40,390.75,145.83,0.0000,-53.190,-22.569,-7.3780,-5.4459,-6.3063,-60.377,0.0000,-101.57,-70.649,-42.682,-62.363
3.000000000000,0.50797E+07,0.50874E+06,0.79242E+06,0.91446E+06,0.93040E+06,0.48589E+06,0.15486E+07,0.21453E+06,0.72564E+06,0.11562E+06,0.29280E+06,0.32093E+06,0.0000,-21247.,-12683.,-2751.8,-4709.6,-9611.5,-38046.,-813.59,-36887.,-10331.,-14171.,-2298.8,12.069,429.96,392.05,160.03,58.139,294.26,337.16,0.0000,1131.4,299.64,673.94,246.33,0.0000,-87.992,-38.585,-11.678,-8.7217,-10.050,-107.36,0.0000,-180.97,-118.95,-83.133,-104.98
4.000000000000,0.37026E+07,0.32180E+06,0.57908E+06,0.69420E+06,0.59228E+06,0.36724E+06,0.12272E+07,0.17957E+06,0.54013E+06,88215.,0.21336E+06,0.24936E+06,0.0000,-21184.,-12417.,-2470.4,-4758.4,-9347.4,-37372.,-803.18,-35346.,-9650.1,-15036.,-2348.0,16.390,583.90,549.44,216.82,78.946,399.49,485.25,0.0000,1613.7,415.74,965.32,341.77,0.0000,-122.92,-54.926,-15.842,-11.964,-13.604,-161.83,0.0000,-284.02,-164.95,-126.60,-145.13
5.000000000000,0.26230E+07,0.23085E+06,0.41825E+06,0.49573E+06,0.40242E+06,0.28302E+06,0.91094E+06,0.14442E+06,0.40719E+06,67720.,0.14902E+06,0.18988E+06,0.0000,-20664.,-12182.,-2274.3,-4801.9,-9122.0,-38401.,-791.41,-34378.,-9075.8,-13784.,-2398.4,20.503,730.42,666.02,270.76,98.749,499.39,627.44,0.0000,2076.2,526.70,1244.9,432.99,0.0000,-156.51,-69.801,-19.801,-15.095,-16.938,-217.90,0.0000,-396.81,-209.38,-171.96,-183.17
6.000000000000,0.19153E+07,0.17236E+06,0.31310E+06,0.37822E+06,0.30067E+06,0.21221E+06,0.69587E+06,0.10948E+06,0.31277E+06,51201.,0.11142E+06,0.14147E+06,0.0000,-20099.,-11935.,-2134.5,-4840.4,-8912.3,-39548.,-778.82,-34770.,-8723.9,-13011.,-2421.2,24.393,868.98,792.37,321.83,117.48,594.00,760.82,0.0000,2510.5,632.85,1507.9,520.25,0.0000,-188.42,-84.091,-23.548,-18.086,-20.068,-265.10,0.0000,-499.21,-251.90,-225.65,-219.40
7.000000000000,0.15076E+07,0.13452E+06,0.25290E+06,0.29703E+06,0.25375E+06,0.16972E+06,0.53501E+06,83547.,0.24621E+06,40997.,90423.,0.11216E+06,0.0000,-19569.,-11700.,-2026.8,-4874.3,-8715.6,-38962.,-766.70,-35489.,-8420.3,-12288.,-2437.9,28.083,1000.5,912.24,370.46,135.25,684.36,891.14,0.0000,2933.7,735.69,1764.5,604.80,0.0000,-218.84,-97.419,-27.108,-20.945,-23.030,-310.51,0.0000,-595.77,-293.09,-279.82,-254.42
8.000000000000,0.12473E+07,0.10877E+06,0.19976E+06,0.23936E+06,0.20912E+06,0.13873E+06,0.43604E+06,70463.,0.20539E+06,32950.,76335.,91448.,0.0000,-19065.,-11478.,-1941.2,-4904.0,-8549.7,-38141.,-755.19,-35521.,-8144.6,-11608.,-2450.3,31.587,1125.3,1026.0,416.80,152.12,770.74,1017.9,0.0000,3344.5,835.68,2014.2,686.99,0.0000,-247.70,-109.80,-30.494,-23.673,-25.840,-354.69,0.0000,-682.67,-333.38,-332.96,-288.44
9.000000000000,0.10894E+07,84569.,0.16692E+06,0.20407E+06,0.16133E+06,0.11296E+06,0.36668E+06,56730.,0.17402E+06,27303.,64258.,76452.,0.0000,-18573.,-11255.,-1873.6,-4929.1,-8395.8,-37548.,-752.22,-34064.,-7895.7,-10981.,-2464.2,267.72,1436.2,1393.0,592.91,303.65,996.96,1150.2,198.41,3898.6,1074.6,2403.1,906.49,0.0000,-279.57,-128.27,-34.168,-27.793,-29.716,-400.77,-9.1369,-772.97,-380.44,-388.64,-339.99
10.00000000000,0.90072E+06,72476.,0.14413E+06,0.17713E+06,0.13819E+06,94565.,0.32116E+06,44893.,0.15242E+06,21879.,54507.,64705.,0.0000,-18136.,-11052.,-1820.4,-4941.8,-8252.9,-36736.,-747.82,-33469.,-7675.2,-10521.,-2514.8,489.08,1862.9,1806.9,682.42,350.78,1131.0,1286.9,509.30,4384.6,1268.8,2719.1,1071.2,0.0000,-316.10,-149.05,-38.454,-31.401,-33.557,-448.41,-23.455,-865.55,-446.02,-443.25,-398.37
11.00000000000,0.73720E+06,68545.,0.13084E+06,0.14841E+06,0.11421E+06,83421.,0.27581E+06,41201.,0.12903E+06,18859.,47778.,56919.,0.0000,-17780.,-10876.,-1778.9,-4931.8,-8117.6,-35919.,-731.62,-32846.,-7489.7,-10244.,-2558.6,43.579,1552.5,1415.6,580.77,235.91,1084.0,1402.9,0.0000,4620.7,1243.4,2831.3,1049.3,0.0000,-345.40,-150.97,-42.124,-33.206,-35.641,-488.81,0.0000,-943.65,-489.12,-482.40,-423.65
12.00000000000,0.61944E+06,63192.,0.11879E+06,0.12978E+06,0.10326E+06,79419.,0.23763E+06,38851.,0.11332E+06,17569.,41894.,50615.,0.0000,-17485.,-10724.,-1746.0,-4919.2,-7983.4,-35145.,-718.14,-32270.,-7322.8,-9748.6,-2571.5,46.681,1663.0,1516.4,620.69,231.74,1154.7,1507.5,0.0000,4960.9,1327.3,3018.0,1098.4,0.0000,-370.84,-161.31,-45.204,-35.454,-38.238,-525.29,0.0000,-1014.2,-529.43,-517.22,-453.61
13.00000000000,0.54870E+06,59440.,99710.,0.11383E+06,96928.,72829.,0.20663E+06,35850.,0.10097E+06,15764.,37758.,44833.,0.0000,-17223.,-10592.,-1720.1,-4905.1,-7852.5,-34392.,-706.74,-31731.,-7172.2,-9275.9,-2581.1,49.527,1764.4,1608.8,661.33,243.63,1231.4,1599.7,0.0000,5268.3,1421.4,3203.7,1173.8,0.0000,-394.15,-170.72,-48.067,-37.648,-40.775,-557.40,0.0000,-1076.5,-568.80,-547.02,-485.35
14.00000000000,0.48982E+06,55267.,87331.,0.10184E+06,90778.,64383.,0.18512E+06,32083.,91325.,14276.,34559.,38148.,0.0000,-17040.,-10478.,-1699.8,-4890.0,-7729.9,-33673.,-696.72,-31224.,-7034.6,-8844.2,-2591.1,52.192,1859.3,1695.4,699.98,254.00,1300.6,1599.7,0.0000,5311.4,1511.1,3227.6,1245.3,0.0000,-415.75,-179.46,-50.769,-39.686,-43.201,-557.41,0.0000,-1078.5,-606.80,-547.56,-515.54
15.00000000000,0.45789E+06,48018.,74126.,92109.,82674.,54157.,0.16376E+06,28205.,80514.,12713.,31628.,34299.,0.0000,-16855.,-10377.,-1681.8,-4874.3,-7615.1,-32992.,-687.63,-30760.,-6908.7,-8458.0,-2601.1,54.700,1948.6,1776.8,736.97,264.99,1367.8,1600.2,0.0000,5354.4,1598.2,3253.0,1315.6,0.0000,-435.99,-187.59,-53.326,-41.604,-45.528,-557.57,0.0000,-1080.7,-643.41,-547.43,-544.55
16.00000000000,0.43595E+06,43363.,69191.,84991.,79108.,48680.,0.14662E+06,22379.,73874.,11596.,29561.,31104.,0.0000,-16684.,-10288.,-1667.6,-4858.4,-7500.8,-32311.,-679.17,-30324.,-6792.8,-8097.4,-2611.4,57.074,2033.2,1854.0,772.36,275.83,1432.8,1604.4,0.0000,5406.3,1682.4,3284.5,1384.0,0.0000,-454.96,-195.20,-55.758,-43.412,-47.761,-559.03,0.0000,-1085.3,-678.69,-547.80,-572.50
17.00000000000,0.42081E+06,38827.,65502.,80157.,75255.,42135.,0.13330E+06,18329.,67643.,10183.,28315.,28353.,0.0000,-16534.,-10209.,-1657.8,-4842.3,-7379.9,-31659.,-671.23,-29928.,-6742.0,-7779.0,-2622.4,59.311,2112.9,1926.6,806.04,286.34,1495.8,1625.6,0.0000,5505.0,1763.7,3345.1,1450.4,0.0000,-472.70,-202.30,-58.060,-45.107,-49.898,-566.42,0.0000,-1100.9,-712.79,-552.65,-599.32
18.00000000000,0.40835E+06,33445.,61660.,74994.,73424.,39102.,0.12380E+06,16705.,61714.,8894.1,26469.,26258.,0.0000,-16403.,-10138.,-1651.6,-4826.0,-7271.5,-31059.,-663.70,-29561.,-6633.6,-7496.6,-2645.2,61.417,2188.0,1995.1,838.03,296.35,1557.7,1686.6,0.0000,5715.5,1843.5,3474.5,1515.8,0.0000,-489.29,-208.92,-60.238,-46.693,-51.938,-587.69,0.0000,-1142.4,-746.34,-568.75,-625.58
19.00000000000,0.39749E+06,30216.,54711.,68951.,69021.,36645.,0.11940E+06,16135.,57280.,8523.7,25014.,25070.,0.0000,-16284.,-10075.,-1647.2,-4809.6,-7172.7,-30516.,-656.51,-29217.,-6563.9,-7241.2,-2664.9,63.419,2259.3,2060.1,868.64,305.98,1614.5,1686.6,0.0000,5750.7,1931.4,3500.6,1587.8,0.0000,-504.95,-215.17,-62.314,-48.190,-53.900,-587.69,0.0000,-1144.2,-783.09,-567.20,-654.54
20.00000000000,0.37773E+06,27796.,51165.,64916.,61176.,33945.,0.11375E+06,15611.,55205.,8282.2,24301.,23754.,0.0000,-16175.,-10018.,-1645.5,-4793.8,-7081.5,-30015.,-649.64,-28887.,-6487.4,-7006.2,-2676.8,65.315,2326.8,2121.7,897.84,315.18,1669.0,1686.6,0.0000,5784.7,2039.4,3532.8,1676.6,0.0000,-519.70,-221.03,-64.288,-49.611,-55.781,-587.69,0.0000,-1146.1,-828.19,-566.47,-690.33
21.00000000000,0.34972E+06,25206.,50248.,61511.,53428.,32245.,0.10788E+06,15166.,53244.,7939.2,23213.,22497.,0.0000,-16073.,-9968.0,-1645.5,-4778.6,-6995.7,-29483.,-643.09,-28582.,-6414.4,-6789.2,-2686.3,67.111,2390.8,2180.0,925.71,323.90,1721.1,1686.6,0.0000,5817.5,2167.5,3571.1,1781.9,0.0000,-533.59,-226.53,-66.164,-50.958,-57.585,-587.69,0.0000,-1148.2,-881.65,-566.46,-732.99
22.00000000000,0.33807E+06,22132.,47827.,58795.,42032.,31736.,0.10429E+06,14933.,49942.,7623.4,21426.,21204.,0.0000,-15977.,-9922.7,-1647.1,-4763.8,-6915.1,-28977.,-636.88,-28312.,-6346.9,-6589.4,-2695.1,68.820,2451.7,2235.5,952.38,332.20,1771.2,1686.6,0.0000,5849.4,2326.1,3618.5,1912.2,0.0000,-546.74,-231.70,-67.955,-52.238,-59.319,-587.69,0.0000,-1149.5,-947.69,-567.48,-786.07
23.00000000000,0.32634E+06,19178.,45456.,56604.,37272.,30326.,0.10092E+06,14471.,46660.,7422.8,19526.,20095.,0.0000,-15887.,-9881.8,-1649.6,-4749.3,-6838.5,-28505.,-630.98,-28059.,-6284.6,-6409.8,-2703.8,70.438,2509.3,2288.1,977.83,340.06,1819.0,1686.6,0.0000,5880.3,2504.3,3671.7,2058.8,0.0000,-559.13,-236.51,-69.658,-53.448,-60.981,-587.69,0.0000,-1150.6,-1022.0,-569.18,-845.96
24.00000000000,0.30273E+06,17861.,37832.,53985.,33732.,27847.,97867.,13967.,44391.,7163.9,17879.,18953.,0.0000,-15806.,-9843.7,-1653.0,-4734.8,-6765.4,-28064.,-625.37,-27820.,-6232.7,-6248.6,-2712.4,71.967,2563.8,2337.7,1002.1,347.49,1864.7,1686.6,0.0000,5909.9,2690.9,3727.4,2212.1,0.0000,-570.77,-240.94,-71.273,-54.585,-62.571,-587.69,0.0000,-1151.5,-1099.8,-571.10,-908.93
25.00000000000,0.27313E+06,15612.,36587.,51164.,30064.,26378.,93448.,13489.,42480.,6744.3,16769.,18024.,0.0000,-15729.,-9807.8,-1656.8,-4720.2,-6695.4,-27631.,-620.00,-27596.,-6191.0,-6100.0,-2721.0,73.413,2615.3,2384.7,1025.2,354.53,1908.5,1686.6,0.0000,5938.3,2879.2,3783.7,2367.0,0.0000,-581.73,-245.05,-72.807,-55.655,-64.096,-587.69,0.0000,-1152.1,-1178.5,-573.10,-972.83
26.00000000000,0.23581E+06,14734.,36308.,48002.,26498.,24729.,89733.,12987.,40247.,6400.3,15126.,17158.,0.0000,-15656.,-9774.0,-1661.2,-4705.6,-6629.3,-27216.,-614.83,-27386.,-6149.3,-5961.9,-2729.5,74.789,2664.3,2429.4,1047.3,361.22,1950.4,1686.6,0.0000,5965.7,3066.0,3839.5,2520.5,0.0000,-592.13,-248.89,-74.272,-56.666,-65.563,-587.69,0.0000,-1152.5,-1257.2,-575.46,-1036.5
27.00000000000,0.20449E+06,14445.,36184.,43486.,24527.,23002.,85348.,12586.,37718.,6311.0,14706.,16409.,0.0000,-15593.,-9742.5,-1666.1,-4690.9,-6566.3,-26827.,-609.87,-27196.,-6110.7,-5834.1,-2738.1,76.103,2711.1,2472.1,1068.5,367.61,1990.8,1686.6,0.0000,5992.1,3249.3,3894.2,2671.1,0.0000,-602.02,-252.54,-75.673,-57.624,-66.977,-587.69,0.0000,-1152.8,-1334.8,-578.02,-1099.3
28.00000000000,0.18187E+06,14444.,32456.,39356.,22948.,22463.,77930.,12179.,35967.,6366.1,13785.,15110.,0.0000,-15532.,-9712.9,-1671.7,-4676.3,-6505.5,-26461.,-605.11,-27020.,-6076.7,-5717.5,-2747.1,77.336,2755.1,2512.2,1088.7,373.62,2029.2,1686.6,0.0000,6017.3,3427.2,3947.4,2817.4,0.0000,-611.25,-255.92,-76.997,-58.517,-68.326,-587.69,0.0000,-1153.0,-1410.5,-580.91,-1160.6
29.00000000000,0.17285E+06,14349.,28798.,36255.,22088.,22271.,71424.,11809.,32407.,6314.8,12459.,14351.,0.0000,-15470.,-9685.0,-1682.3,-4661.9,-6446.9,-26118.,-600.52,-26858.,-6047.9,-5609.2,-2756.4,78.499,2796.5,2549.9,1107.9,379.29,2065.9,1686.6,0.0000,6041.3,3599.1,3998.7,2958.8,0.0000,-619.89,-259.06,-78.251,-59.352,-69.617,-587.69,0.0000,-1153.0,-1484.2,-584.05,-1220.2
30.00000000000,0.15317E+06,13903.,28684.,33328.,20167.,21805.,65867.,11510.,31043.,6111.8,11612.,13545.,0.0000,-15408.,-9658.6,-1691.0,-4647.7,-6390.5,-25794.,-596.10,-26703.,-6023.7,-5508.5,-2765.8,79.644,2837.3,2587.1,1126.7,384.87,2102.0,1686.6,0.0000,6065.0,3767.4,4049.0,3097.1,0.0000,-628.35,-262.11,-79.484,-60.169,-70.888,-587.69,0.0000,-1153.0,-1556.7,-587.56,-1279.8
31.00000000000,0.12879E+06,13504.,28722.,31322.,18851.,21702.,61825.,11441.,29305.,6086.5,10920.,12920.,0.0000,-15346.,-9633.5,-1698.7,-4633.7,-6336.3,-25490.,-591.80,-26557.,-6003.3,-5414.7,-2775.2,80.772,2877.4,2623.8,1145.3,390.36,2137.4,1686.6,0.0000,6088.2,3932.4,4098.3,3232.7,0.0000,-636.66,-265.08,-80.699,-60.969,-72.141,-587.69,0.0000,-1153.0,-1628.2,-591.80,-1339.0
32.00000000000,0.11703E+06,13456.,24879.,29323.,17548.,20363.,55896.,10851.,27552.,5797.3,10210.,12177.,0.0000,-15286.,-9609.7,-1706.1,-4620.0,-6284.2,-25203.,-587.63,-26418.,-5986.6,-5327.4,-2784.7,81.832,2915.2,2658.2,1162.9,395.53,2171.3,1686.6,0.0000,6110.4,4091.9,4145.9,3363.9,0.0000,-644.40,-267.81,-81.847,-61.716,-73.340,-587.69,0.0000,-1152.9,-1697.8,-596.24,-1396.7
33.00000000000,0.11262E+06,13466.,21625.,25890.,16218.,19909.,50222.,10371.,26263.,5651.4,9444.1,11399.,0.0000,-15226.,-9587.9,-1713.5,-4606.5,-6234.5,-24933.,-583.57,-26286.,-5982.4,-5246.1,-2794.0,82.827,2950.7,2690.5,1179.6,400.38,2203.5,1686.6,0.0000,6131.3,4220.3,4184.3,3469.5,0.0000,-651.60,-270.33,-82.931,-62.410,-74.486,-587.69,0.0000,-1152.6,-1754.4,-601.95,-1444.1
34.00000000000,0.10216E+06,13398.,21570.,24168.,15925.,18634.,48345.,9845.5,25220.,5605.9,8456.1,10656.,0.0000,-15168.,-9568.2,-1721.0,-4593.3,-6186.9,-24686.,-579.63,-26170.,-5981.1,-5170.3,-2802.6,83.764,2984.1,2721.0,1195.6,404.96,2234.3,1686.6,0.0000,6149.8,4220.3,4184.3,3469.5,0.0000,-658.34,-272.66,-83.958,-63.059,-75.584,-587.69,0.0000,-1150.8,-1757.4,-602.26,-1447.4
35.00000000000,93188.,13085.,21520.,22857.,15934.,17578.,44073.,9236.9,24050.,5519.9,7961.1,9891.4,0.0000,-15111.,-9549.9,-1728.6,-4580.3,-6141.6,-24452.,-575.80,-26058.,-5974.8,-5099.3,-2810.7,84.657,3015.9,2750.0,1210.9,409.32,2264.0,1686.6,0.0000,6167.7,4220.5,4184.3,3469.6,0.0000,-664.72,-274.84,-84.940,-63.673,-76.645,-587.69,0.0000,-1149.0,-1760.5,-602.62,-1450.5
36.00000000000,85037.,13008.,18320.,21722.,15852.,16268.,40857.,8533.0,23353.,5413.0,7482.1,8763.4,0.0000,-15055.,-9532.8,-1736.5,-4567.6,-6098.8,-24230.,-572.07,-25950.,-5977.4,-5033.0,-2818.5,85.488,3045.5,2777.0,1225.3,413.38,2292.1,1686.6,0.0000,6184.6,4221.0,4184.5,3470.0,0.0000,-670.61,-276.80,-85.861,-64.238,-77.655,-587.69,0.0000,-1147.3,-1763.4,-603.04,-1453.4
37.00000000000,81008.,13020.,14464.,19607.,15688.,13945.,38660.,8080.8,21931.,5169.2,7229.8,8531.3,0.0000,-15001.,-9516.6,-1744.4,-4555.1,-6057.7,-24021.,-568.44,-25847.,-5974.4,-4972.4,-2826.0,86.284,3073.8,2802.8,1239.2,417.27,2319.4,1686.6,0.0000,6201.1,4223.6,4185.3,3472.2,0.0000,-676.22,-278.63,-86.747,-64.775,-78.635,-587.69,0.0000,-1145.8,-1767.1,-603.60,-1456.7
38.00000000000,77535.,12470.,14366.,18109.,15643.,12629.,35138.,7346.7,20611.,4953.0,7026.7,8367.1,0.0000,-14947.,-9501.1,-1752.5,-4542.8,-6018.0,-23828.,-564.92,-25747.,-5968.3,-4918.4,-2833.3,87.026,3100.3,2826.9,1252.4,420.90,2345.3,1686.6,0.0000,6216.8,4235.8,4188.9,3482.2,0.0000,-681.49,-280.28,-87.581,-65.271,-79.572,-587.69,0.0000,-1144.4,-1774.6,-604.66,-1463.2
39.00000000000,73309.,11996.,14393.,17654.,15613.,12118.,32382.,6726.2,19622.,4937.9,6936.9,8233.8,0.0000,-14896.,-9486.9,-1760.8,-4530.8,-5979.6,-23654.,-561.50,-25651.,-5993.3,-4869.0,-2840.3,87.741,3125.7,2850.1,1265.2,424.40,2370.4,1686.6,0.0000,6232.2,4256.2,4195.0,3499.0,0.0000,-686.53,-281.82,-88.385,-65.746,-80.483,-587.69,0.0000,-1143.1,-1784.7,-606.18,-1472.8
40.00000000000,69686.,11973.,14452.,17043.,15620.,11815.,30481.,5618.7,18595.,4805.6,6814.6,7846.3,0.0000,-14849.,-9473.2,-1769.1,-4519.0,-5942.5,-23495.,-558.15,-25559.,-5993.0,-4824.9,-2846.9,88.432,3150.3,2872.6,1277.6,427.79,2394.9,1686.6,0.0000,6248.0,4350.0,4223.0,3576.0,0.0000,-691.37,-283.28,-89.165,-66.201,-81.373,-587.69,0.0000,-1142.8,-1825.5,-611.31,-1508.4
41.00000000000,68529.,11952.,14494.,15604.,15550.,11167.,28538.,4649.7,18483.,4621.9,6895.6,7251.7,0.0000,-14804.,-9459.7,-1777.5,-4507.5,-5906.6,-23344.,-554.89,-25470.,-5992.4,-4786.3,-2853.3,89.085,3173.6,2893.8,1289.6,430.99,2418.5,1686.6,0.0000,6263.4,4449.7,4252.8,3658.0,0.0000,-695.92,-284.61,-89.909,-66.628,-82.234,-587.69,0.0000,-1142.7,-1869.0,-617.48,-1546.7
42.00000000000,67875.,11887.,14371.,15010.,15548.,10088.,26482.,4199.3,18311.,4479.1,6832.6,7016.2,0.0000,-14759.,-9446.5,-1786.0,-4496.2,-5871.9,-23200.,-551.68,-25385.,-5992.2,-4750.1,-2859.4,89.698,3195.4,2913.7,1300.9,434.00,2440.9,1686.6,0.0000,6276.9,4449.7,4252.8,3658.0,0.0000,-700.15,-285.81,-90.610,-67.025,-83.056,-587.69,0.0000,-1141.4,-1870.5,-619.75,-1550.2
43.00000000000,67716.,11859.,14304.,14456.,15554.,9270.9,24941.,3647.7,17411.,4394.7,6795.7,6834.1,0.0000,-14714.,-9433.5,-1794.5,-4485.2,-5839.8,-23063.,-548.52,-25304.,-5992.4,-4715.7,-2865.1,90.278,3216.1,2932.6,1311.7,436.84,2462.5,1686.6,0.0000,6289.9,4449.7,4252.8,3658.0,0.0000,-704.13,-286.90,-91.279,-67.398,-83.850,-587.69,0.0000,-1140.3,-1871.9,-621.98,-1553.3
44.00000000000,67239.,11846.,14276.,14131.,15560.,8805.5,23965.,3328.6,16921.,4175.6,6795.6,6668.7,0.0000,-14670.,-9421.2,-1803.1,-4474.3,-5809.1,-22933.,-545.43,-25225.,-5993.4,-4683.2,-2870.5,90.863,3237.0,2951.6,1322.5,439.72,2484.1,1686.6,0.0000,6302.9,4449.7,4252.8,3658.0,0.0000,-708.17,-288.01,-91.951,-67.774,-84.644,-587.69,0.0000,-1139.2,-1873.6,-624.17,-1556.3
45.00000000000,67122.,11713.,14205.,13805.,15490.,8748.6,22893.,3217.7,16511.,4092.8,6794.9,6466.7,0.0000,-14627.,-9409.4,-1811.7,-4463.7,-5779.1,-22809.,-542.40,-25150.,-5994.7,-4652.4,-2875.4,91.424,3256.9,2969.8,1333.0,442.47,2504.9,1686.6,0.0000,6315.5,4449.7,4252.8,3658.0,0.0000,-712.00,-289.04,-92.597,-68.131,-85.415,-587.69,0.0000,-1138.2,-1875.2,-626.32,-1559.0
46.00000000000,66941.,11711.,14152.,13569.,15432.,8687.1,22250.,3114.6,16290.,4083.8,6793.5,6246.7,0.0000,-14584.,-9398.1,-1820.5,-4453.4,-5750.0,-22691.,-539.43,-25076.,-5995.7,-4623.2,-2880.1,91.948,3275.6,2986.8,1343.0,445.04,2524.9,1686.6,0.0000,6327.5,4449.7,4252.8,3658.0,0.0000,-715.53,-289.95,-93.208,-68.462,-86.159,-587.69,0.0000,-1137.3,-1876.6,-628.43,-1561.5
47.00000000000,66803.,11552.,14160.,13323.,15402.,8132.6,21486.,3080.4,15162.,4050.1,6791.4,6214.8,0.0000,-14542.,-9387.0,-1829.2,-4443.2,-5722.2,-22578.,-536.51,-25005.,-5996.6,-4595.5,-2884.4,92.466,3294.1,3003.6,1352.8,447.59,2544.6,1686.6,0.0000,6339.4,4449.7,4252.8,3658.0,0.0000,-719.01,-290.83,-93.811,-68.789,-86.892,-587.69,0.0000,-1136.4,-1877.9,-630.59,-1563.9
48.00000000000,66725.,11458.,14071.,13314.,15401.,8123.1,20685.,3048.3,14825.,4037.2,6789.0,6210.3,0.0000,-14501.,-9376.0,-1838.1,-4433.2,-5696.0,-22470.,-533.65,-24936.,-5997.1,-4569.4,-2888.4,92.950,3311.3,3019.3,1362.1,449.97,2563.4,1686.6,0.0000,6350.7,4449.7,4252.8,3658.0,0.0000,-722.20,-291.60,-94.379,-69.090,-87.597,-587.69,0.0000,-1135.6,-1879.0,-633.20,-1566.0
49.00000000000,66536.,11433.,14007.,13255.,15326.,8133.6,20559.,3036.4,14842.,4028.1,6785.9,6177.5,0.0000,-14459.,-9365.3,-1846.9,-4423.5,-5672.5,-22368.,-530.86,-24870.,-5997.5,-4544.6,-2892.2,93.377,3326.5,3033.2,1370.7,452.08,2580.8,1686.6,0.0000,6361.2,4449.7,4252.8,3658.0,0.0000,-724.93,-292.18,-94.891,-69.350,-88.317,-587.69,0.0000,-1134.8,-1880.1,-636.29,-1568.0
50.00000000000,66398.,11362.,14008.,13212.,15332.,8111.4,20450.,2987.3,14873.,4025.4,6782.8,6175.5,0.0000,-14418.,-9354.7,-1855.8,-4413.9,-5653.0,-22269.,-528.15,-24805.,-5999.0,-4521.1,-2895.6,93.759,3340.1,3045.6,1378.7,453.97,2597.2,1686.6,0.0000,6371.1,4449.7,4252.8,3658.0,0.0000,-727.30,-292.62,-95.360,-69.577,-89.005,-587.69,0.0000,-1134.1,-1880.9,-639.35,-1569.8
51.00000000000,66375.,11274.,13960.,13187.,15337.,8085.1,20010.,2966.1,14888.,4022.1,6779.3,6157.7,0.0000,-14377.,-9344.2,-1864.8,-4404.6,-5635.1,-22175.,-525.50,-24742.,-6007.2,-4498.9,-2898.8,94.142,3353.7,3058.1,1386.6,455.86,2613.5,1686.6,0.0000,6380.9,4449.7,4252.8,3658.0,0.0000,-729.63,-293.05,-95.828,-69.804,-89.625,-587.69,0.0000,-1133.4,-1881.5,-642.62,-1571.5
52.00000000000,66346.,11189.,13953.,13209.,15263.,8101.4,19852.,2955.4,14829.,4003.7,6826.4,6157.9,0.0000,-14337.,-9334.0,-1873.8,-4395.4,-5617.3,-22086.,-523.06,-24680.,-6012.2,-4478.0,-2901.9,94.544,3368.1,3071.1,1395.1,457.85,2631.0,1686.6,0.0000,6391.5,4449.7,4252.8,3658.0,0.0000,-732.10,-293.56,-96.326,-70.047,-90.280,-587.69,0.0000,-1132.8,-1882.0,-646.09,-1573.1
53.00000000000,66296.,11187.,13969.,13212.,15177.,8092.9,19764.,2928.6,14402.,3993.3,6824.8,6171.3,0.0000,-14297.,-9323.9,-1882.8,-4386.5,-5599.6,-22000.,-520.50,-24620.,-6015.8,-4458.3,-2905.0,94.891,3380.5,3082.4,1402.5,459.57,2646.3,1686.6,0.0000,6400.7,4449.7,4252.8,3658.0,0.0000,-734.14,-293.96,-96.758,-70.250,-90.850,-587.69,0.0000,-1132.2,-1882.4,-649.49,-1574.5
54.00000000000,66298.,11202.,13996.,13139.,15063.,8076.9,19738.,2916.0,14413.,3985.0,6803.5,6173.7,0.0000,-14258.,-9313.9,-1891.9,-4377.7,-5581.9,-21917.,-517.97,-24562.,-6018.8,-4444.8,-2907.9,95.218,3392.1,3093.0,1409.5,461.20,2661.0,1686.6,0.0000,6409.6,4449.7,4252.8,3658.0,0.0000,-736.01,-294.29,-97.167,-70.438,-91.396,-587.69,0.0000,-1131.6,-1882.8,-652.80,-1575.8
55.00000000000,66226.,11215.,13977.,13136.,15048.,8111.3,19697.,2916.7,14418.,3985.0,6798.1,6142.2,0.0000,-14219.,-9304.0,-1901.0,-4369.1,-5564.6,-21838.,-515.50,-24505.,-6021.3,-4433.2,-2910.6,95.526,3403.1,3103.0,1416.4,462.73,2675.2,1686.6,0.0000,6418.2,4449.7,4252.8,3658.0,0.0000,-737.74,-294.57,-97.559,-70.614,-91.926,-587.69,0.0000,-1131.1,-1883.0,-656.23,-1577.0
56.00000000000,66161.,11229.,13937.,13037.,14721.,8065.3,19704.,2890.7,14397.,3967.6,6777.1,6124.6,0.0000,-14181.,-9294.4,-1910.2,-4360.6,-5547.9,-21763.,-513.23,-24449.,-6023.8,-4420.5,-2913.1,95.881,3415.7,3114.5,1423.8,464.48,2690.5,1686.6,0.0000,6427.4,4449.7,4252.8,3658.0,0.0000,-739.81,-294.99,-97.995,-70.824,-92.490,-587.69,0.0000,-1130.6,-1883.2,-659.57,-1578.1
57.00000000000,66132.,11250.,13965.,13041.,14598.,8065.0,19705.,2874.8,14346.,3963.6,6759.6,6123.5,0.0000,-14145.,-9285.0,-1919.4,-4352.3,-5531.3,-21690.,-510.86,-24395.,-6026.3,-4407.7,-2915.5,96.202,3427.2,3125.0,1430.7,466.07,2704.8,1686.6,0.0000,6436.1,4449.7,4252.8,3658.0,0.0000,-741.63,-295.31,-98.397,-71.011,-93.021,-587.69,0.0000,-1130.1,-1883.4,-662.83,-1579.1
58.00000000000,66032.,11251.,13987.,12901.,14356.,8075.4,19636.,2859.5,14289.,3957.2,6749.2,6125.6,0.0000,-14113.,-9275.8,-1928.4,-4344.2,-5518.3,-21621.,-508.51,-24342.,-6033.5,-4395.4,-2917.6,96.480,3437.0,3134.0,1437.0,467.46,2718.1,1686.6,0.0000,6444.1,4449.7,4252.8,3658.0,0.0000,-743.11,-295.50,-98.756,-71.166,-93.423,-587.69,0.0000,-1129.7,-1883.2,-666.00,-1580.0
59.00000000000,65960.,11213.,13961.,12868.,14244.,8055.5,19638.,2859.9,14279.,3953.2,6746.0,6131.2,0.0000,-14081.,-9266.7,-1936.4,-4336.2,-5517.6,-21554.,-506.21,-24291.,-6042.6,-4383.8,-2919.5,96.752,3446.7,3142.9,1443.2,468.81,2731.2,1686.6,0.0000,6452.0,4449.7,4252.8,3658.0,0.0000,-744.55,-295.68,-99.109,-71.318,-93.789,-587.69,0.0000,-1129.3,-1882.9,-669.09,-1580.8
60.00000000000,65910.,11178.,13973.,12797.,14187.,8030.2,19569.,2860.6,14287.,3947.7,6740.1,6130.3,0.0000,-14049.,-9257.8,-1943.3,-4328.3,-5520.0,-21490.,-503.95,-24240.,-6049.0,-4372.7,-2921.3,97.006,3455.8,3151.1,1449.2,470.08,2743.8,1686.6,0.0000,6459.6,4449.7,4252.8,3658.0,0.0000,-745.84,-295.81,-99.443,-71.456,-94.128,-587.69,0.0000,-1128.9,-1882.5,-672.09,-1581.8
61.00000000000,65533.,11109.,13897.,12779.,14148.,7991.3,19576.,2838.0,14295.,3945.8,6723.0,6129.5,0.0000,-14017.,-9249.0,-1949.3,-4320.5,-5521.9,-21430.,-501.73,-24191.,-6054.3,-4362.2,-2924.4,97.230,3463.7,3158.4,1454.7,471.20,2755.7,1686.6,0.0000,6466.8,4449.7,4252.8,3658.0,0.0000,-746.90,-295.84,-99.747,-71.574,-94.434,-587.69,0.0000,-1128.5,-1882.1,-675.02,-1582.6
62.00000000000,65454.,11082.,13906.,12786.,14107.,7938.4,19581.,2825.9,14250.,3938.9,6748.4,6121.6,0.0000,-13985.,-9240.3,-1954.7,-4312.8,-5522.9,-21372.,-499.54,-24143.,-6059.2,-4352.2,-2937.8,97.436,3471.1,3165.1,1460.0,472.24,2767.1,1686.6,0.0000,6473.7,4449.7,4252.8,3658.0,0.0000,-747.83,-295.83,-100.04,-71.679,-94.722,-587.69,0.0000,-1128.2,-1881.7,-677.88,-1583.0
63.00000000000,65248.,11092.,13829.,12776.,13983.,7940.9,19587.,2826.7,14147.,3939.8,6729.0,6097.0,0.0000,-13952.,-9231.7,-1959.6,-4305.2,-5523.4,-21318.,-497.38,-24096.,-6064.0,-4342.7,-2945.4,97.595,3476.8,3170.2,1464.6,473.05,2777.4,1686.6,0.0000,6479.9,4449.7,4252.8,3658.0,0.0000,-748.40,-295.68,-100.28,-71.750,-94.965,-587.69,0.0000,-1127.8,-1881.2,-680.68,-1583.3
64.00000000000,64931.,11096.,13785.,12631.,13986.,7916.9,19559.,2821.3,14075.,3934.3,6729.2,6092.3,0.0000,-13921.,-9223.2,-1964.1,-4297.7,-5523.4,-21268.,-495.25,-24050.,-6068.6,-4334.4,-2950.1,97.719,3481.2,3174.3,1468.8,473.69,2786.7,1686.6,0.0000,6485.6,4449.7,4252.8,3658.0,0.0000,-748.73,-295.42,-100.48,-71.796,-95.175,-587.69,0.0000,-1127.5,-1881.0,-683.31,-1583.6
65.00000000000,64825.,11046.,13755.,12598.,13988.,7865.5,19483.,2808.5,14033.,3926.1,6737.5,6092.2,0.0000,-13891.,-9214.7,-1968.3,-4290.3,-5523.0,-21219.,-493.14,-24005.,-6073.1,-4345.0,-2954.1,97.883,3487.0,3179.6,1473.4,474.52,2797.0,1686.6,0.0000,6491.7,4449.7,4252.8,3658.0,0.0000,-749.39,-295.28,-100.72,-71.872,-95.413,-587.69,0.0000,-1127.2,-1880.8,-685.52,-1583.8
66.00000000000,64632.,10944.,13528.,12527.,13928.,7817.8,19412.,2806.3,14003.,3918.6,6695.2,6092.1,0.0000,-13861.,-9206.3,-1972.1,-4282.9,-5522.3,-21172.,-491.05,-23961.,-6077.6,-4341.1,-2958.5,98.031,3492.3,3184.4,1477.8,475.28,2806.7,1686.6,0.0000,6497.6,4449.7,4252.8,3658.0,0.0000,-749.92,-295.10,-100.95,-71.937,-95.635,-587.69,0.0000,-1126.9,-1880.5,-687.66,-1583.9
67.00000000000,64377.,10897.,13438.,12605.,13870.,7748.4,19319.,2806.9,14025.,3919.1,6664.2,6092.2,0.0000,-13831.,-9198.0,-1975.8,-4275.7,-5521.3,-21126.,-488.98,-23918.,-6082.0,-4338.2,-2962.7,98.145,3496.4,3188.1,1481.8,475.87,2815.7,1686.6,0.0000,6503.1,4449.7,4252.8,3658.0,0.0000,-750.20,-294.82,-101.15,-71.978,-95.828,-587.69,0.0000,-1126.6,-1880.2,-689.74,-1583.9
68.00000000000,64216.,10851.,13382.,12612.,13848.,7752.1,19298.,2797.2,14033.,3912.1,6654.2,6092.4,0.0000,-13801.,-9189.8,-1979.2,-4268.5,-5520.1,-21081.,-486.93,-23876.,-6086.5,-4335.8,-2966.4,98.211,3498.7,3190.3,1485.1,476.23,2823.5,1686.6,0.0000,6507.8,4449.7,4252.8,3658.0,0.0000,-750.10,-294.40,-101.29,-71.984,-95.979,-587.69,0.0000,-1126.3,-1879.9,-691.75,-1583.8
69.00000000000,64127.,10791.,13337.,12619.,13794.,7762.0,19235.,2790.1,14040.,3905.2,6646.2,6092.7,0.0000,-13772.,-9181.6,-1982.5,-4261.5,-5518.7,-21038.,-485.24,-23835.,-6091.1,-4333.7,-2969.9,99.011,3514.6,3204.7,1491.2,478.37,2834.3,1686.6,0.0000,6514.3,4449.7,4252.8,3658.0,0.0000,-752.88,-295.11,-101.73,-72.268,-96.233,-587.69,0.0000,-1126.1,-1879.5,-693.71,-1583.7
70.00000000000,63927.,10732.,13282.,12619.,13696.,7764.4,18983.,2790.7,13999.,3899.1,6612.9,6092.9,0.0000,-13742.,-9173.8,-1985.7,-4254.5,-5517.1,-20996.,-483.18,-23793.,-6095.6,-4332.1,-2972.8,98.777,3518.9,3208.6,1495.1,479.00,2843.2,1686.6,0.0000,6519.7,4449.7,4252.8,3658.0,0.0000,-753.17,-294.87,-101.93,-72.317,-96.421,-587.69,0.0000,-1125.9,-1879.1,-695.62,-1583.5
71.00000000000,63824.,10739.,13258.,12527.,13587.,7708.2,18799.,2791.3,13890.,3889.0,6598.7,6075.7,0.0000,-13713.,-9166.0,-1988.7,-4247.6,-5515.4,-20955.,-481.11,-23753.,-6100.3,-4330.9,-2975.4,98.871,3522.2,3211.7,1498.7,479.49,2851.4,1686.6,0.0000,6524.6,4449.7,4252.8,3658.0,0.0000,-753.23,-294.53,-102.10,-72.347,-96.584,-587.69,0.0000,-1125.7,-1878.7,-697.49,-1583.2
72.00000000000,63762.,10745.,13179.,12477.,13576.,7728.1,18777.,2791.9,13846.,3878.4,6588.6,6075.7,0.0000,-13683.,-9158.3,-1991.6,-4240.7,-5513.9,-20916.,-479.08,-23714.,-6105.2,-4329.8,-2977.8,98.931,3524.4,3213.6,1501.8,479.82,2858.8,1686.6,0.0000,6529.1,4449.7,4252.8,3658.0,0.0000,-753.04,-294.10,-102.23,-72.352,-96.720,-587.69,0.0000,-1125.4,-1878.2,-699.30,-1582.9
73.00000000000,63606.,10679.,13031.,12397.,13508.,7742.4,18659.,2787.5,13767.,3871.9,6570.6,6076.0,0.0000,-13653.,-9150.6,-1994.4,-4233.9,-5512.7,-20878.,-477.11,-23675.,-6110.1,-4328.9,-2980.1,98.961,3525.4,3214.6,1504.4,480.00,2865.3,1686.6,0.0000,6533.1,4449.7,4252.8,3658.0,0.0000,-752.63,-293.58,-102.34,-72.334,-96.827,-587.69,0.0000,-1125.2,-1877.7,-701.08,-1582.5
74.00000000000,62401.,10647.,13034.,12383.,12917.,7750.9,18484.,2760.4,13697.,3847.6,6565.7,6067.7,0.0000,-13623.,-9142.9,-1997.1,-4227.2,-5511.5,-20840.,-475.17,-23637.,-6114.8,-4328.1,-2982.2,98.971,3525.8,3214.9,1506.8,480.09,2871.3,1686.6,0.0000,6536.7,4449.7,4252.8,3658.0,0.0000,-752.14,-293.00,-102.43,-72.304,-96.917,-587.69,0.0000,-1125.0,-1877.1,-702.99,-1582.1
75.00000000000,62244.,10592.,13038.,12334.,12196.,7764.7,18476.,2758.1,13702.,3821.2,6564.0,6058.3,0.0000,-13592.,-9135.1,-1999.7,-4220.5,-5510.0,-20804.,-473.27,-23600.,-6119.5,-4330.3,-2984.1,98.954,3525.2,3214.4,1508.7,480.04,2876.6,1686.6,0.0000,6539.9,4449.7,4252.8,3658.0,0.0000,-751.43,-292.34,-102.48,-72.253,-96.981,-587.69,0.0000,-1124.8,-1876.6,-704.76,-1581.7
76.00000000000,62045.,10465.,13042.,12301.,12198.,7782.3,18381.,2743.9,13626.,3794.4,6545.8,6058.9,0.0000,-13562.,-9127.3,-2002.2,-4213.8,-5508.4,-20769.,-471.38,-23563.,-6124.1,-4336.1,-2985.9,98.918,3523.9,3213.2,1510.5,479.91,2881.4,1686.6,0.0000,6542.9,4449.7,4252.8,3658.0,0.0000,-750.57,-291.62,-102.52,-72.190,-97.031,-587.69,0.0000,-1124.6,-1876.0,-706.36,-1581.2
77.00000000000,61874.,10340.,13044.,12257.,12200.,7788.9,18341.,2736.6,13626.,3784.9,6527.4,6057.1,0.0000,-13532.,-9119.5,-2004.6,-4207.2,-5506.5,-20735.,-469.52,-23528.,-6128.7,-4343.3,-2987.6,98.893,3523.0,3212.4,1512.3,479.82,2886.4,1686.6,0.0000,6545.9,4449.7,4252.8,3658.0,0.0000,-749.79,-290.93,-102.57,-72.134,-97.085,-587.69,0.0000,-1124.4,-1875.4,-707.78,-1580.7
78.00000000000,61810.,10167.,13041.,12150.,12167.,7794.9,18345.,2734.8,13622.,3779.0,6512.3,6047.3,0.0000,-13502.,-9111.7,-2006.9,-4200.7,-5504.5,-20701.,-467.67,-23492.,-6133.2,-4349.4,-2989.1,98.865,3522.0,3211.5,1514.0,479.73,2891.3,1686.6,0.0000,6548.9,4449.7,4252.8,3658.0,0.0000,-748.99,-290.24,-102.62,-72.078,-97.136,-587.69,0.0000,-1124.2,-1874.9,-709.09,-1580.3
79.00000000000,61876.,10074.,12962.,12013.,12065.,7798.2,18350.,2723.5,13567.,3774.9,6500.8,6012.4,0.0000,-13472.,-9103.9,-2009.2,-4194.2,-5502.4,-20669.,-465.84,-23458.,-6137.7,-4359.0,-2991.4,98.837,3521.0,3210.6,1515.7,479.63,2896.0,1686.6,0.0000,6551.8,4449.7,4252.8,3658.0,0.0000,-748.19,-289.54,-102.66,-72.021,-97.184,-587.69,0.0000,-1124.0,-1874.2,-710.14,-1579.7
80.00000000000,61876.,9989.5,12929.,12014.,12054.,7742.8,18354.,2703.5,13505.,3766.4,6485.4,5997.2,0.0000,-13442.,-9096.1,-2011.4,-4187.7,-5500.1,-20637.,-464.03,-23425.,-6142.1,-4367.4,-2995.5,98.803,3519.8,3209.5,1517.3,479.50,2900.6,1686.6,0.0000,6554.5,4449.7,4252.8,3658.0,0.0000,-747.33,-288.83,-102.70,-71.960,-97.224,-587.69,0.0000,-1123.8,-1873.6,-711.15,-1579.1
81.00000000000,61751.,9895.3,12814.,11952.,12056.,7749.0,18359.,2682.4,13440.,3760.2,6479.6,5992.9,0.0000,-13412.,-9088.3,-2013.5,-4181.3,-5497.7,-20606.,-462.24,-23392.,-6146.5,-4373.2,-2998.5,98.746,3517.8,3207.6,1518.6,479.26,2904.5,1686.6,0.0000,6556.9,4449.7,4252.8,3658.0,0.0000,-746.27,-288.06,-102.71,-71.884,-97.244,-587.69,0.0000,-1123.6,-1873.0,-712.12,-1578.4
82.00000000000,61551.,9805.6,12689.,11953.,11980.,7754.8,18363.,2681.1,13418.,3753.5,6467.9,5973.0,0.0000,-13383.,-9080.6,-2015.6,-4174.9,-5495.3,-20576.,-460.59,-23360.,-6150.9,-4378.1,-3000.6,98.864,3522.0,3211.5,1522.5,479.99,2913.3,1686.6,0.0000,6562.3,4449.7,4252.8,3658.0,0.0000,-746.52,-287.79,-102.91,-71.936,-97.432,-587.69,0.0000,-1123.5,-1872.6,-713.05,-1577.8
83.00000000000,61331.,9800.7,12641.,11957.,11917.,7698.6,18368.,2664.4,13421.,3747.9,6453.0,5962.7,0.0000,-13353.,-9072.8,-2017.7,-4168.6,-5492.8,-20547.,-458.81,-23328.,-6155.2,-4382.6,-3002.2,98.816,3520.3,3209.9,1523.8,479.67,2917.2,1686.6,0.0000,6564.7,4449.7,4252.8,3658.0,0.0000,-745.52,-287.04,-102.93,-71.866,-97.455,-587.69,0.0000,-1123.4,-1872.2,-713.95,-1577.1
84.00000000000,61067.,9728.7,12616.,11923.,11911.,7682.3,18372.,2645.8,13331.,3737.7,6436.2,5961.6,0.0000,-13324.,-9065.1,-2019.7,-4162.3,-5490.1,-20518.,-457.02,-23296.,-6159.5,-4386.9,-3003.4,98.841,3521.2,3210.7,1526.1,479.82,2922.9,1686.6,0.0000,6568.1,4449.7,4252.8,3658.0,0.0000,-745.06,-286.51,-103.02,-71.850,-97.536,-587.69,0.0000,-1123.2,-1871.8,-714.81,-1576.4
85.00000000000,60927.,9611.9,12577.,11874.,11913.,7619.5,18254.,2631.5,13299.,3728.5,6418.3,5926.4,0.0000,-13295.,-9057.6,-2021.7,-4156.1,-5487.4,-20490.,-455.26,-23265.,-6163.7,-4391.1,-3004.6,98.860,3521.8,3211.3,1528.2,479.94,2928.3,1686.6,0.0000,6571.4,4449.7,4252.8,3658.0,0.0000,-744.56,-285.96,-103.10,-71.831,-97.610,-587.69,0.0000,-1123.1,-1871.3,-715.65,-1575.7
86.00000000000,60912.,9524.1,12563.,11782.,11915.,7570.7,18145.,2617.1,13246.,3684.0,6417.5,5891.4,0.0000,-13266.,-9050.2,-2023.6,-4149.9,-5484.5,-20463.,-453.52,-23235.,-6167.9,-4395.1,-3005.6,98.855,3521.6,3211.2,1530.1,479.95,2933.1,1686.6,0.0000,6574.3,4449.7,4252.8,3658.0,0.0000,-743.88,-285.35,-103.16,-71.795,-97.664,-587.69,0.0000,-1123.0,-1870.8,-716.46,-1575.0
87.00000000000,60839.,9492.0,12509.,11741.,11917.,7472.8,18149.,2607.1,13224.,3668.7,6416.7,5890.3,0.0000,-13238.,-9042.8,-2025.5,-4143.8,-5481.6,-20437.,-451.81,-23205.,-6171.9,-4399.0,-3006.5,98.797,3519.6,3209.3,1531.2,479.70,2936.6,1686.6,0.0000,6576.5,4449.7,4252.8,3658.0,0.0000,-742.80,-284.58,-103.17,-71.720,-97.673,-587.69,0.0000,-1122.8,-1870.3,-717.25,-1574.3
88.00000000000,59747.,9387.1,12400.,11745.,11919.,7473.1,18153.,2593.5,13212.,3647.3,6392.3,5822.9,0.0000,-13209.,-9035.4,-2027.4,-4137.7,-5478.5,-20411.,-450.12,-23175.,-6176.0,-4402.8,-3007.3,98.698,3516.1,3206.1,1531.7,479.26,2939.1,1686.6,0.0000,6578.0,4449.7,4252.8,3658.0,0.0000,-741.41,-283.70,-103.14,-71.616,-97.647,-587.69,0.0000,-1122.7,-1869.8,-718.02,-1573.6
89.00000000000,59416.,9233.8,12257.,11724.,11920.,7478.0,18092.,2593.9,13168.,3625.9,6386.3,5775.7,0.0000,-13180.,-9028.0,-2029.2,-4131.7,-5475.4,-20385.,-448.46,-23145.,-6179.9,-4406.5,-3008.0,98.593,3512.3,3202.7,1532.1,478.79,2941.3,1686.6,0.0000,6579.3,4449.7,4252.8,3658.0,0.0000,-739.99,-282.80,-103.10,-71.509,-97.612,-587.69,0.0000,-1122.5,-1869.2,-718.77,-1573.0
90.00000000000,59381.,9172.3,12162.,11590.,11922.,7482.5,18025.,2580.4,13149.,3615.1,6385.6,5755.8,0.0000,-13152.,-9020.5,-2030.9,-4125.6,-5472.1,-20360.,-446.83,-23116.,-6183.8,-4410.1,-3008.7,98.457,3507.5,3198.2,1532.0,478.16,2942.6,1686.6,0.0000,6580.2,4449.7,4252.8,3658.0,0.0000,-738.30,-281.82,-103.02,-71.378,-97.551,-587.69,0.0000,-1122.3,-1868.7,-719.49,-1572.5
91.00000000000,59380.,9152.8,12114.,11593.,11868.,7486.6,17941.,2576.6,13112.,3609.9,6385.0,5714.7,0.0000,-13123.,-9013.0,-2032.6,-4119.6,-5468.8,-20336.,-445.22,-23088.,-6187.6,-4413.6,-3009.2,98.327,3502.9,3194.0,1531.9,477.56,2943.9,1686.6,0.0000,6581.0,4449.7,4252.8,3658.0,0.0000,-736.66,-280.85,-102.96,-71.252,-97.487,-587.69,0.0000,-1122.2,-1868.1,-720.20,-1572.0
92.00000000000,59380.,9016.1,12085.,11596.,11820.,7500.3,17945.,2561.4,12997.,3595.0,6384.2,5682.1,0.0000,-13094.,-9005.5,-2034.2,-4113.6,-5466.6,-20312.,-443.64,-23060.,-6191.4,-4417.0,-3009.7,98.202,3498.4,3190.0,1532.0,476.99,2945.4,1686.6,0.0000,6581.9,4449.7,4252.8,3658.0,0.0000,-735.06,-279.90,-102.89,-71.130,-97.431,-587.69,0.0000,-1122.0,-1867.4,-720.89,-1571.4
93.00000000000,59364.,8995.9,11749.,11571.,11522.,7511.2,17834.,2555.5,12982.,3586.9,6365.2,5673.2,0.0000,-13066.,-8998.2,-2035.8,-4107.7,-5464.9,-20289.,-442.59,-23032.,-6195.3,-4420.4,-3010.6,98.731,3512.5,3203.0,1539.9,479.36,2961.6,1686.6,0.33393E-01,6591.7,4449.7,4252.9,3658.0,0.0000,-737.35,-280.44,-103.37,-71.389,-97.870,-587.69,-0.15366E-02,-1122.1,-1866.9,-721.56,-1570.9
94.00000000000,59299.,8971.5,11689.,11498.,11274.,7516.5,17767.,2555.3,12985.,3584.2,6349.9,5656.9,0.0000,-13038.,-8991.1,-2037.4,-4101.9,-5462.7,-20266.,-440.95,-23004.,-6199.0,-4423.7,-3010.9,98.595,3512.4,3202.7,1541.4,478.95,2965.6,1686.6,0.0000,6594.1,4449.7,4252.8,3658.0,0.0000,-736.68,-279.85,-103.42,-71.355,-97.903,-587.69,0.0000,-1122.0,-1866.3,-722.22,-1570.3
95.00000000000,59197.,8811.1,11691.,11462.,11209.,7476.2,17722.,2555.6,12952.,3581.3,6317.5,5641.3,0.0000,-13010.,-8984.2,-2039.0,-4096.1,-5460.2,-20244.,-439.25,-22977.,-6202.6,-4426.9,-3011.0,98.524,3509.9,3200.4,1542.1,478.64,2968.0,1686.6,0.0000,6595.6,4449.7,4252.8,3658.0,0.0000,-735.50,-279.07,-103.40,-71.274,-97.880,-587.69,0.0000,-1121.9,-1865.8,-722.86,-1569.8
96.00000000000,59042.,8689.8,11591.,11343.,11129.,7471.7,17650.,2571.7,12895.,3559.7,6294.3,5632.1,0.0000,-12982.,-8977.2,-2040.6,-4090.3,-5457.7,-20222.,-437.59,-22951.,-6206.1,-4430.1,-3011.0,98.429,3506.5,3197.3,1542.4,478.21,2969.8,1686.6,0.0000,6596.7,4449.7,4252.8,3658.0,0.0000,-734.13,-278.23,-103.36,-71.176,-97.836,-587.69,0.0000,-1121.7,-1865.2,-723.49,-1569.3
97.00000000000,58748.,8603.2,11520.,11329.,11130.,7475.8,17584.,2553.5,12782.,3553.4,6285.3,5557.5,0.0000,-12954.,-8970.1,-2042.1,-4084.6,-5454.9,-20200.,-435.99,-22925.,-6209.5,-4433.2,-3011.1,98.280,3501.2,3192.5,1541.9,477.52,2970.3,1686.6,0.0000,6597.0,4449.7,4252.8,3658.0,0.0000,-732.37,-277.24,-103.27,-71.039,-97.748,-587.69,0.0000,-1121.6,-1864.7,-724.10,-1568.7
98.00000000000,58586.,8427.4,11466.,11255.,11079.,7479.2,17482.,2547.6,12679.,3544.5,6284.7,5540.7,0.0000,-12925.,-8963.0,-2043.5,-4078.8,-5452.0,-20179.,-434.43,-22899.,-6213.0,-4436.1,-3014.6,98.108,3495.0,3186.9,1541.1,476.71,2970.1,1686.6,0.0000,6597.0,4449.7,4252.8,3658.0,0.0000,-730.43,-276.18,-103.16,-70.885,-97.638,-587.69,0.0000,-1121.4,-1864.1,-724.70,-1568.0
99.00000000000,58552.,8338.5,11411.,11243.,10784.,7455.3,17444.,2520.6,12616.,3552.3,6266.1,5513.6,0.0000,-12896.,-8955.8,-2045.0,-4073.1,-5449.0,-20159.,-432.91,-22874.,-6216.4,-4438.8,-3018.4,97.917,3488.2,3180.7,1540.0,475.82,2969.4,1686.6,0.0000,6596.6,4449.7,4252.8,3658.0,0.0000,-728.35,-275.08,-103.02,-70.718,-97.512,-587.69,0.0000,-1121.3,-1863.5,-725.28,-1567.3
100.0000000000,57678.,8321.8,11392.,11200.,9910.0,7414.8,17447.,2513.3,12531.,3548.1,6245.3,5505.8,0.0000,-12867.,-8948.7,-2046.3,-4067.4,-5445.9,-20138.,-431.41,-22849.,-6219.7,-4441.2,-3021.1,97.762,3482.7,3175.6,1539.3,475.09,2969.5,1686.6,0.0000,6596.7,4449.7,4252.8,3658.0,0.0000,-726.54,-274.07,-102.92,-70.577,-97.413,-587.69,0.0000,-1121.2,-1862.8,-725.86,-1566.6
101.0000000000,57389.,8194.7,11332.,11105.,9882.8,7306.9,17411.,2506.8,12391.,3535.1,6227.7,5477.9,0.0000,-12838.,-8941.5,-2047.6,-4061.7,-5442.7,-20119.,-429.94,-22825.,-6223.1,-4443.7,-3023.2,97.665,3479.3,3172.5,1539.5,474.65,2971.0,1686.6,0.0000,6597.6,4449.7,4252.8,3658.0,0.0000,-725.16,-273.24,-102.87,-70.478,-97.359,-587.69,0.0000,-1121.0,-1862.2,-726.42,-1566.0
102.0000000000,57389.,8131.1,11127.,11046.,9883.7,7262.9,17298.,2495.8,12328.,3516.3,6225.0,5473.9,0.0000,-12809.,-8934.4,-2048.8,-4056.1,-5439.4,-20099.,-428.50,-22803.,-6226.2,-4446.0,-3027.5,97.540,3474.8,3168.4,1539.2,474.07,2971.7,1686.6,0.0000,6598.1,4449.7,4252.8,3658.0,0.0000,-723.57,-272.32,-102.80,-70.359,-97.282,-587.69,0.0000,-1120.9,-1861.5,-726.97,-1565.2
103.0000000000,57358.,8043.9,11075.,10935.,9880.7,7113.2,17249.,2493.3,12329.,3512.4,6224.5,5457.5,0.0000,-12781.,-8927.3,-2049.9,-4050.4,-5436.0,-20080.,-427.09,-22782.,-6229.2,-4448.3,-3033.1,97.392,3469.5,3163.6,1538.6,473.39,2971.9,1686.6,0.0000,6598.2,4449.7,4252.8,3658.0,0.0000,-721.81,-271.35,-102.71,-70.224,-97.186,-587.69,0.0000,-1120.8,-1860.9,-727.51,-1564.4
104.0000000000,57323.,7947.7,11073.,10803.,9610.0,7002.3,17140.,2464.1,12298.,3507.9,6206.9,5416.1,0.0000,-12752.,-8920.2,-2051.1,-4044.8,-5432.6,-20061.,-425.70,-22766.,-6232.2,-4450.6,-3037.3,97.235,3464.0,3158.5,1537.9,472.65,2971.8,1686.6,0.0000,6598.2,4449.7,4252.8,3658.0,0.0000,-719.98,-270.35,-102.60,-70.082,-97.078,-587.69,0.0000,-1120.7,-1860.1,-728.04,-1563.5
105.0000000000,57297.,7906.5,11070.,10789.,9561.2,6888.5,17073.,2453.8,12261.,3492.7,6159.6,5348.2,0.0000,-12723.,-8913.1,-2052.1,-4039.2,-5429.2,-20043.,-424.34,-22754.,-6236.1,-4452.8,-3045.9,97.018,3456.2,3151.5,1536.3,471.63,2970.1,1686.6,0.0000,6597.2,4449.7,4252.8,3658.0,0.0000,-717.71,-269.19,-102.43,-69.897,-96.918,-587.69,0.0000,-1120.4,-1859.3,-728.56,-1562.7
106.0000000000,57147.,7690.9,11003.,10702.,9561.9,6772.3,16944.,2441.4,12262.,3483.2,6144.6,5349.1,0.0000,-12694.,-8905.9,-2053.1,-4033.6,-5425.6,-20025.,-423.00,-22742.,-6240.2,-4455.0,-3062.6,96.786,3448.0,3144.0,1534.5,470.53,2968.0,1686.6,0.0000,6596.0,4449.7,4252.8,3658.0,0.0000,-715.34,-267.99,-102.25,-69.702,-96.744,-587.69,0.0000,-1120.2,-1858.5,-729.06,-1561.9
107.0000000000,56982.,7622.7,10992.,10684.,9528.1,6763.0,16759.,2425.8,12273.,3483.4,6126.0,5347.6,0.0000,-12665.,-8898.7,-2054.1,-4028.0,-5422.0,-20007.,-421.67,-22731.,-6244.0,-4457.1,-3071.9,96.553,3439.6,3136.4,1532.7,469.43,2965.9,1686.6,0.0000,6594.7,4449.7,4252.8,3658.0,0.0000,-712.95,-266.78,-102.07,-69.506,-96.566,-587.69,0.0000,-1119.9,-1857.7,-729.55,-1561.1
108.0000000000,56768.,7557.4,10947.,10608.,9476.7,6695.8,16707.,2426.0,12198.,3479.8,6081.6,5320.5,0.0000,-12636.,-8891.5,-2054.9,-4022.4,-5418.2,-19989.,-420.61,-22719.,-6247.6,-4459.2,-3079.6,96.619,3442.0,3138.5,1535.1,469.78,2971.4,1686.6,0.0000,6598.1,4449.7,4252.8,3658.0,0.0000,-712.78,-266.41,-102.19,-69.526,-96.638,-587.69,0.0000,-1119.7,-1856.9,-730.03,-1560.3
109.0000000000,56628.,7520.7,10919.,10589.,9477.6,6615.2,16696.,2424.1,12144.,3475.2,6069.5,5315.6,0.0000,-12608.,-8884.5,-2055.8,-4016.9,-5414.3,-19972.,-419.26,-22708.,-6250.9,-4461.2,-3086.5,96.506,3438.0,3134.9,1534.9,469.25,2972.1,1686.6,0.0000,6598.5,4449.7,4252.8,3658.0,0.0000,-711.29,-265.55,-102.12,-69.417,-96.550,-587.69,0.0000,-1119.4,-1856.2,-730.49,-1559.5
110.0000000000,56222.,7439.1,10880.,10576.,9411.8,6626.4,16602.,2404.0,12145.,3450.1,6069.1,5307.4,0.0000,-12579.,-8877.6,-2056.6,-4011.4,-5410.4,-19955.,-417.90,-22699.,-6254.0,-4463.2,-3092.9,96.381,3433.5,3130.8,1534.5,468.67,2972.5,1686.6,0.0000,6598.8,4449.7,4252.8,3658.0,0.0000,-709.71,-264.66,-102.04,-69.300,-96.449,-587.69,0.0000,-1119.1,-1855.4,-730.95,-1558.7
111.0000000000,55356.,7209.5,10778.,10577.,9297.6,6627.9,16457.,2382.3,12134.,3427.8,6019.4,5267.4,0.0000,-12551.,-8870.7,-2057.4,-4005.9,-5406.4,-19938.,-416.57,-22689.,-6257.0,-4465.1,-3099.0,96.220,3427.8,3125.6,1533.6,467.92,2972.1,1686.6,0.0000,6598.5,4449.7,4252.8,3658.0,0.0000,-707.87,-263.67,-101.93,-69.157,-96.317,-587.69,0.0000,-1118.9,-1854.7,-731.39,-1557.9
112.0000000000,55304.,7132.9,10707.,10579.,9237.5,6628.8,16328.,2363.7,12059.,3414.0,5954.8,5244.4,0.0000,-12523.,-8863.7,-2058.1,-4000.4,-5402.4,-19922.,-415.27,-22679.,-6259.9,-4467.0,-3104.9,96.035,3421.2,3119.6,1532.4,467.05,2971.0,1686.6,0.0000,6597.9,4449.7,4252.8,3658.0,0.0000,-705.87,-262.63,-101.79,-68.998,-96.163,-587.69,0.0000,-1118.6,-1853.9,-731.82,-1557.2
113.0000000000,55136.,6939.9,10574.,10579.,9187.1,6629.4,16331.,2332.3,12060.,3405.0,5934.2,5244.2,0.0000,-12495.,-8856.7,-2058.8,-3994.9,-5398.2,-19906.,-414.00,-22668.,-6262.8,-4468.9,-3110.6,95.820,3413.5,3112.6,1530.7,466.04,2969.1,1686.6,0.0000,6596.8,4449.7,4252.8,3658.0,0.0000,-703.64,-261.50,-101.63,-68.817,-95.981,-587.69,0.0000,-1118.3,-1853.1,-732.24,-1556.6
114.0000000000,54905.,6900.4,10408.,10541.,9158.2,6633.3,16332.,2316.7,12069.,3380.2,5929.3,5226.5,0.0000,-12468.,-8849.8,-2059.4,-3989.4,-5393.9,-19890.,-412.75,-22658.,-6265.6,-4470.7,-3116.1,95.691,3408.9,3108.4,1530.3,465.43,2969.3,1686.6,0.0000,6597.0,4449.7,4252.8,3658.0,0.0000,-702.05,-260.61,-101.54,-68.697,-95.866,-587.69,0.0000,-1118.0,-1852.4,-732.65,-1556.0
115.0000000000,54738.,6803.2,10383.,10442.,9150.8,6638.9,16272.,2281.1,12070.,3366.3,5914.3,5225.9,0.0000,-12440.,-8842.8,-2059.9,-3984.0,-5389.6,-19874.,-411.53,-22647.,-6268.4,-4472.5,-3121.5,95.578,3404.9,3104.7,1530.0,464.91,2969.9,1686.6,0.0000,6597.4,4449.7,4252.8,3658.0,0.0000,-700.58,-259.77,-101.48,-68.590,-95.762,-587.69,0.0000,-1117.7,-1851.6,-733.06,-1555.4
116.0000000000,54737.,6660.8,10278.,10353.,9009.5,6640.2,16154.,2272.9,12070.,3365.3,5896.2,5203.6,0.0000,-12412.,-8835.9,-2060.4,-3978.6,-5385.2,-19858.,-410.31,-22637.,-6271.1,-4474.3,-3126.6,95.416,3399.1,3099.5,1529.0,464.15,2969.3,1686.6,0.0000,6597.0,4449.7,4252.8,3658.0,0.0000,-698.75,-258.80,-101.36,-68.447,-95.615,-587.69,0.0000,-1117.4,-1850.8,-733.45,-1554.7
117.0000000000,54666.,6597.6,10243.,10353.,8848.9,6641.1,16005.,2258.6,12019.,3361.5,5894.7,5191.5,0.0000,-12385.,-8829.0,-2060.9,-3973.2,-5380.7,-19843.,-409.10,-22626.,-6273.7,-4476.0,-3131.6,95.206,3391.6,3092.6,1527.4,463.16,2967.4,1686.6,0.0000,6595.9,4449.7,4252.8,3658.0,0.0000,-696.58,-257.70,-101.20,-68.270,-95.426,-587.69,0.0000,-1117.1,-1850.0,-733.84,-1554.1
118.0000000000,54495.,6564.7,10210.,10354.,8815.8,6627.9,15929.,2246.7,11929.,3358.9,5894.3,5184.3,0.0000,-12359.,-8822.6,-2061.3,-3967.9,-5376.3,-19828.,-408.62,-22616.,-6276.8,-4477.7,-3137.2,97.371,3445.3,3143.1,1549.8,471.22,3008.5,1686.6,0.0000,6620.4,4449.7,4252.8,3658.0,0.0000,-706.82,-261.26,-102.72,-69.317,-96.642,-587.69,0.0000,-1117.3,-1849.3,-734.22,-1553.5
119.0000000000,54021.,6496.3,10144.,10359.,8792.4,6577.6,15932.,2219.9,11922.,3353.5,5888.1,5162.0,0.0000,-12336.,-8817.8,-2062.1,-3962.9,-5371.9,-19813.,-408.61,-22605.,-6280.1,-4479.3,-3143.4,136.84,3616.9,3501.9,1598.7,495.78,3097.7,1686.6,0.31823,6669.2,4450.0,4253.2,3658.4,0.0000,-723.05,-273.00,-105.27,-71.023,-99.217,-587.69,-0.14628E-01,-1118.0,-1848.5,-734.59,-1553.0
120.0000000000,53258.,6396.2,10178.,10372.,8716.0,6581.8,15935.,2214.4,11872.,3348.5,5853.2,5130.5,0.0000,-12317.,-8814.6,-2063.3,-3958.2,-5368.0,-19798.,-406.97,-22595.,-6282.6,-4480.9,-3147.7,99.655,3550.1,3237.1,1595.4,510.21,3093.8,1686.6,0.0000,6671.9,4449.7,4252.8,3658.0,0.0000,-727.41,-268.32,-105.81,-71.591,-99.198,-587.69,0.0000,-1117.8,-1847.8,-734.96,-1552.3
121.0000000000,52952.,6340.8,10200.,10388.,8703.6,6589.1,15876.,2212.8,11878.,3343.4,5830.0,5110.6,0.0000,-12298.,-8811.5,-2064.4,-3953.6,-5364.4,-19784.,-405.26,-22585.,-6284.8,-4482.5,-3151.5,99.706,3552.0,3238.8,1596.0,487.78,3094.7,1686.6,0.0000,6672.4,4449.7,4252.8,3658.0,0.0000,-727.28,-268.04,-105.86,-71.443,-99.098,-587.69,0.0000,-1117.5,-1847.1,-735.32,-1551.7
122.0000000000,52875.,6161.5,10169.,10370.,8708.1,6602.1,15794.,2191.0,11889.,3320.6,5808.0,5087.0,0.0000,-12281.,-8808.6,-2065.7,-3949.0,-5360.9,-19770.,-404.19,-22575.,-6287.2,-4484.1,-3155.8,335.68,3782.4,3416.9,1629.3,491.26,3113.6,1686.6,2.8038,6689.2,4449.7,4252.8,3658.0,0.0000,-736.12,-273.87,-106.87,-72.280,-99.500,-587.69,-0.12887,-1117.4,-1846.3,-735.67,-1551.0
123.0000000000,52646.,6139.2,10122.,10186.,8634.0,6612.6,15565.,2175.1,11897.,3310.3,5791.6,5075.7,0.0000,-12264.,-8806.2,-2067.0,-3944.4,-5357.0,-19756.,-402.72,-22565.,-6289.5,-4485.6,-3159.7,101.37,3611.4,3293.0,1611.4,493.35,3116.1,1686.6,0.0000,6685.1,4449.7,4252.8,3658.0,0.0000,-738.52,-271.76,-107.24,-72.590,-99.528,-587.69,0.0000,-1117.2,-1845.6,-736.02,-1550.4
124.0000000000,51380.,6102.5,10114.,10048.,8519.4,6623.0,15546.,2174.6,11872.,3301.1,5779.5,5063.4,0.0000,-12249.,-8803.8,-2068.3,-3939.9,-5353.0,-19742.,-401.32,-22556.,-6291.6,-4487.1,-3163.4,101.48,3615.0,3296.3,1613.1,493.53,3119.3,1686.6,0.0000,6687.0,4449.7,4252.8,3658.0,0.0000,-738.81,-271.66,-107.35,-72.644,-99.497,-587.69,0.0000,-1116.9,-1844.9,-736.36,-1549.7
125.0000000000,51287.,6047.9,10019.,9843.8,8398.2,6634.8,15421.,2154.3,11820.,3297.1,5764.8,5019.0,0.0000,-12233.,-8801.1,-2069.6,-3935.3,-5348.8,-19728.,-400.02,-22546.,-6293.9,-4488.6,-3167.0,101.41,3612.8,3294.3,1613.4,493.14,3120.9,1686.6,0.0000,6688.0,4449.7,4252.8,3658.0,0.0000,-737.92,-271.13,-107.33,-72.581,-99.411,-587.69,0.0000,-1116.7,-1844.1,-736.69,-1549.1
126.0000000000,51199.,5928.1,9969.7,9759.7,8394.5,6647.8,15290.,2132.1,11644.,3297.8,5742.0,4977.1,0.0000,-12216.,-8798.1,-2070.6,-3930.7,-5344.3,-19715.,-398.79,-22536.,-6296.1,-4490.0,-3170.7,101.26,3607.4,3289.4,1613.0,492.42,3121.4,1686.6,0.0000,6688.3,4449.7,4252.8,3658.0,0.0000,-736.38,-270.36,-107.24,-72.454,-99.291,-587.69,0.0000,-1116.4,-1843.4,-737.03,-1548.7
127.0000000000,51141.,5838.7,9924.8,9572.3,8372.7,6640.3,15190.,2117.1,11642.,3298.5,5722.1,4932.2,0.0000,-12199.,-8794.8,-2071.5,-3926.0,-5339.8,-19702.,-397.60,-22526.,-6298.3,-4491.5,-3174.3,101.06,3600.2,3282.8,1612.0,491.48,3121.1,1686.6,0.0000,6688.2,4449.7,4252.8,3658.0,0.0000,-734.46,-269.46,-107.10,-72.289,-99.146,-587.69,0.0000,-1116.1,-1842.6,-737.35,-1548.2
128.0000000000,51117.,5692.0,9616.2,9534.1,8282.2,6556.3,15178.,2103.8,11580.,3293.0,5701.6,4923.1,0.0000,-12181.,-8791.2,-2072.3,-3921.3,-5335.0,-19688.,-396.45,-22516.,-6300.6,-4492.9,-3177.9,100.82,3591.7,3275.0,1610.6,490.35,3120.2,1686.6,0.0000,6687.7,4449.7,4252.8,3658.0,0.0000,-732.26,-268.44,-106.93,-72.097,-98.980,-587.69,0.0000,-1115.8,-1841.8,-737.67,-1547.6
129.0000000000,51001.,5524.6,9551.3,9536.1,8226.2,6487.6,15116.,2103.9,11582.,3288.0,5683.6,4923.7,0.0000,-12162.,-8787.4,-2072.9,-3916.6,-5330.1,-19676.,-395.32,-22506.,-6302.9,-4494.3,-3181.4,100.56,3582.3,3266.4,1608.9,489.11,3118.8,1686.6,0.0000,6686.9,4449.7,4252.8,3658.0,0.0000,-729.88,-267.36,-106.74,-71.887,-98.798,-587.69,0.0000,-1115.5,-1841.1,-737.99,-1547.1
130.0000000000,50943.,5392.8,9284.3,9423.1,8168.2,6490.7,14954.,2104.1,11585.,3280.7,5683.3,4916.7,0.0000,-12143.,-8783.4,-2073.5,-3911.9,-5325.2,-19663.,-394.40,-22497.,-6305.3,-4495.6,-3185.1,165.42,3602.6,3322.8,1612.8,494.87,3125.0,1686.6,0.0000,6690.6,4449.7,4252.8,3658.0,0.0000,-731.97,-268.88,-107.05,-72.146,-98.857,-587.69,0.0000,-1115.3,-1840.3,-738.30,-1546.6
131.0000000000,50870.,5389.8,9194.6,9397.1,8139.7,6481.0,14913.,2104.2,11552.,3267.6,5654.9,4895.7,0.0000,-12125.,-8779.9,-2074.1,-3907.3,-5320.1,-19651.,-393.51,-22487.,-6307.7,-4497.0,-3188.7,178.13,3685.5,3382.0,1632.2,505.75,3147.1,1686.6,0.0000,6699.7,4449.7,4252.8,3658.0,0.0000,-735.67,-270.86,-107.61,-72.580,-99.259,-587.69,0.0000,-1115.2,-1839.6,-738.60,-1546.1
132.0000000000,50825.,5384.1,9093.6,9335.8,8047.1,6427.5,14915.,2094.5,11491.,3245.0,5607.6,4887.5,0.0000,-12108.,-8776.6,-2074.7,-3902.7,-5315.1,-19638.,-392.32,-22477.,-6310.0,-4498.3,-3191.8,101.43,3613.5,3295.0,1621.0,493.35,3140.3,1686.6,0.0000,6699.8,4449.7,4252.8,3658.0,0.0000,-734.90,-268.60,-107.60,-72.455,-99.073,-587.69,0.0000,-1114.9,-1838.8,-738.90,-1545.6
133.0000000000,50823.,5278.8,9013.0,9179.3,7906.6,6420.3,14918.,2068.7,11450.,3224.7,5607.4,4840.0,0.0000,-12091.,-8773.1,-2075.3,-3898.2,-5310.0,-19626.,-391.13,-22467.,-6312.3,-4499.6,-3194.8,101.31,3609.2,3291.0,1620.4,492.78,3140.1,1686.6,0.0000,6699.7,4449.7,4252.8,3658.0,0.0000,-733.57,-267.92,-107.52,-72.348,-99.176,-587.69,0.0000,-1114.6,-1838.0,-739.20,-1545.0
134.0000000000,50732.,5177.4,8933.6,9134.5,7907.1,6410.6,14920.,2068.8,11438.,3211.1,5598.4,4821.6,0.0000,-12073.,-8769.4,-2075.8,-3893.6,-5305.0,-19615.,-389.97,-22458.,-6314.5,-4500.9,-3197.8,101.12,3602.2,3284.7,1619.2,491.86,3139.0,1686.6,0.0000,6699.1,4449.7,4252.8,3658.0,0.0000,-731.70,-267.04,-107.38,-72.188,-99.244,-587.69,0.0000,-1114.3,-1837.2,-739.49,-1544.5
135.0000000000,49716.,5171.6,8881.6,9064.7,7893.2,6282.2,14922.,2058.1,11400.,3200.3,5588.0,4773.8,0.0000,-12055.,-8765.5,-2076.3,-3889.1,-5299.8,-19603.,-389.15,-22448.,-6316.9,-4502.2,-3201.0,101.32,3635.1,3336.4,1633.0,501.79,3159.3,1686.6,2.5557,6709.9,4451.9,4254.6,3659.7,0.0000,-732.80,-268.17,-107.67,-72.379,-99.801,-587.69,-0.11741,-1114.3,-1836.4,-739.79,-1544.1
136.0000000000,49779.,5110.0,8842.6,9063.3,7343.2,6255.7,14809.,2041.1,11371.,3196.9,5574.0,4732.6,0.0000,-12037.,-8761.5,-2076.8,-3884.5,-5294.5,-19592.,-388.00,-22438.,-6319.2,-4503.4,-3203.9,101.06,3600.1,3282.7,1622.6,491.65,3148.7,1686.6,0.0000,6704.9,4449.7,4252.8,3658.0,0.0000,-730.37,-266.15,-107.46,-72.105,-99.758,-587.69,0.0000,-1114.0,-1835.6,-740.07,-1543.4
137.0000000000,49474.,5089.6,8760.4,9017.9,6801.0,6213.3,14663.,2019.7,11302.,3192.1,5568.4,4725.7,0.0000,-12019.,-8757.2,-2077.2,-3879.9,-5289.3,-19581.,-386.84,-22429.,-6321.3,-4504.6,-3206.6,100.73,3588.3,3272.0,1619.7,490.08,3144.8,1686.6,0.0000,6702.7,4449.7,4252.8,3658.0,0.0000,-727.52,-264.91,-107.19,-71.847,-99.728,-587.69,0.0000,-1113.8,-1834.8,-740.34,-1542.8
138.0000000000,48446.,5033.5,8658.0,8878.3,6726.1,6215.9,14651.,2001.0,11176.,3183.3,5508.9,4722.0,0.0000,-12000.,-8752.5,-2077.5,-3875.3,-5283.9,-19570.,-385.71,-22419.,-6323.5,-4505.8,-3209.3,100.37,3575.8,3260.5,1616.5,488.41,3140.5,1686.6,0.0000,6700.1,4449.7,4252.8,3658.0,0.0000,-724.51,-263.60,-106.90,-71.574,-99.682,-587.69,0.0000,-1113.6,-1834.0,-740.62,-1542.3
139.0000000000,48288.,4988.4,8621.8,8762.0,6677.7,6217.1,14542.,1980.6,11156.,3175.5,5478.9,4672.5,0.0000,-11980.,-8747.6,-2077.5,-3870.7,-5278.4,-19559.,-384.61,-22409.,-6325.6,-4507.0,-3212.0,100.03,3563.7,3249.5,1613.5,486.79,3136.5,1686.6,0.0000,6697.8,4449.7,4252.8,3658.0,0.0000,-721.58,-262.32,-106.63,-71.309,-99.643,-587.69,0.0000,-1113.3,-1833.2,-740.89,-1541.7
140.0000000000,48217.,4867.9,8615.7,8629.8,6526.9,6191.3,14454.,1976.1,11157.,3175.8,5411.7,4634.3,0.0000,-11961.,-8742.4,-2077.4,-3866.0,-5272.8,-19548.,-383.54,-22400.,-6327.7,-4508.2,-3214.7,99.679,3551.0,3237.9,1610.2,485.11,3132.1,1686.6,0.0000,6695.2,4449.7,4252.8,3658.0,0.0000,-718.53,-261.00,-106.33,-71.033,-99.587,-587.69,0.0000,-1113.1,-1832.4,-741.16,-1541.0
141.0000000000,47935.,4832.3,8607.5,8596.1,6413.7,6127.5,14423.,1958.3,11148.,3171.7,5343.2,4613.6,0.0000,-11940.,-8736.9,-2077.3,-3861.3,-5267.0,-19537.,-382.48,-22390.,-6329.8,-4509.3,-3217.3,99.320,3538.2,3226.3,1606.9,483.40,3127.6,1686.6,0.0000,6692.5,4449.7,4252.8,3658.0,0.0000,-715.45,-259.66,-106.03,-70.754,-99.522,-587.69,0.0000,-1112.9,-1831.5,-741.43,-1540.4
142.0000000000,47912.,4824.1,8599.2,8595.1,6240.9,6047.7,14281.,1958.4,11053.,3169.4,5342.1,4567.6,0.0000,-11919.,-8731.3,-2077.1,-3856.6,-5261.2,-19526.,-381.43,-22381.,-6331.8,-4510.4,-3219.8,98.994,3526.6,3215.7,1604.1,481.86,3123.8,1686.6,0.0000,6690.2,4449.7,4252.8,3658.0,0.0000,-712.60,-258.40,-105.77,-70.499,-99.478,-587.69,0.0000,-1112.7,-1830.7,-741.69,-1539.7
143.0000000000,46948.,4816.4,8562.1,8581.3,6153.0,6046.5,14137.,1958.5,11007.,3149.9,5327.6,4521.4,0.0000,-11898.,-8725.5,-2076.8,-3851.9,-5255.3,-19515.,-380.39,-22371.,-6333.9,-4511.6,-3222.2,98.660,3514.7,3204.8,1601.0,480.27,3119.7,1686.6,0.0000,6687.8,4449.7,4252.8,3658.0,0.0000,-709.69,-257.12,-105.49,-70.238,-99.421,-587.69,0.0000,-1112.4,-1829.8,-741.95,-1539.0
144.0000000000,46702.,4815.3,8520.6,8500.9,6113.7,6046.0,13989.,1954.4,11007.,3141.7,5302.6,4509.6,0.0000,-11878.,-8719.8,-2076.6,-3847.2,-5249.3,-19503.,-379.98,-22361.,-6336.2,-4512.7,-3225.3,128.38,3580.9,3264.4,1627.0,496.29,3160.2,1686.6,10.342,6712.5,4454.8,4257.0,3662.1,0.0000,-714.51,-259.38,-106.38,-70.823,-100.58,-587.69,-0.47496,-1112.6,-1829.0,-742.22,-1538.8
145.0000000000,46561.,4766.5,8526.0,8414.4,6078.2,6049.5,13815.,1940.8,11007.,3139.3,5266.6,4475.4,0.0000,-11858.,-8714.7,-2076.5,-3842.7,-5243.4,-19492.,-378.90,-22352.,-6338.2,-4513.7,-3227.7,99.458,3543.1,3230.8,1617.3,484.22,3153.0,1686.6,0.0000,6707.9,4449.7,4252.8,3658.0,0.0000,-714.45,-258.42,-106.46,-70.764,-100.66,-587.69,0.0000,-1112.4,-1828.2,-742.45,-1537.7
146.0000000000,45792.,4707.1,8542.2,8332.7,6030.7,6054.8,13721.,1940.9,10941.,3128.8,5229.9,4425.7,0.0000,-11840.,-8710.4,-2076.5,-3838.4,-5237.7,-19481.,-378.80,-22342.,-6340.6,-4514.8,-3230.9,307.14,3816.4,3461.9,1671.3,525.79,3219.8,1686.6,142.70,6751.8,4468.5,4269.9,3674.9,0.0000,-730.05,-267.12,-108.42,-72.517,-102.23,-587.69,-6.5531,-1112.6,-1827.4,-742.78,-1538.7
147.0000000000,44807.,4737.5,8571.3,8339.6,5986.0,6063.6,13649.,1925.9,10941.,3113.0,5192.0,4419.7,0.0000,-11826.,-8707.4,-2076.9,-3834.3,-5232.2,-19470.,-377.46,-22333.,-6342.4,-4515.9,-3233.0,102.20,3640.9,3319.9,1645.3,497.44,3194.4,1686.6,0.0000,6732.7,4452.5,4255.6,3663.0,0.0000,-733.31,-264.87,-108.82,-72.689,-102.13,-587.69,0.0000,-1112.5,-1826.6,-742.96,-1536.9
148.0000000000,44673.,4735.7,8587.0,8278.2,5911.2,6072.2,13573.,1923.3,10916.,3107.6,5171.2,4405.6,0.0000,-11812.,-8704.7,-2077.2,-3830.2,-5226.8,-19459.,-376.09,-22324.,-6344.0,-4516.9,-3234.8,102.17,3639.7,3318.8,1643.6,497.10,3190.6,1686.6,0.0000,6730.2,4450.0,4253.2,3658.8,0.0000,-732.66,-264.46,-108.75,-72.649,-102.09,-587.69,0.0000,-1112.3,-1825.7,-743.19,-1535.8
149.0000000000,44320.,4740.3,8575.1,8217.0,5912.8,6077.5,13507.,1923.4,10850.,3108.4,5150.6,4403.0,0.0000,-11797.,-8701.6,-2077.6,-3826.1,-5221.4,-19448.,-374.98,-22315.,-6345.7,-4517.9,-3236.7,102.18,3640.2,3319.3,1644.3,497.18,3192.3,1686.6,11.043,6731.2,4452.4,4252.8,3658.1,0.0000,-732.38,-264.18,-108.78,-72.643,-102.22,-587.69,-0.50707,-1112.1,-1824.9,-743.42,-1535.0
150.0000000000,43844.,4742.3,8526.7,8221.2,5859.6,6081.1,13405.,1923.4,10669.,3095.8,5121.8,4375.2,0.0000,-11783.,-8698.2,-2077.9,-3821.9,-5215.8,-19437.,-373.82,-22306.,-6347.4,-4519.0,-3238.6,101.91,3630.6,3310.5,1641.4,495.90,3187.8,1686.6,0.0000,6728.6,4449.7,4252.8,3658.0,0.0000,-730.06,-263.17,-108.55,-72.435,-102.16,-587.69,0.0000,-1111.9,-1824.0,-743.66,-1534.2
151.0000000000,41848.,4729.9,8488.8,8223.0,5438.1,6033.7,13316.,1907.5,10591.,3085.2,5072.3,4315.6,0.0000,-11767.,-8694.4,-2078.1,-3817.6,-5210.0,-19426.,-372.72,-22297.,-6349.0,-4520.0,-3240.5,101.59,3619.1,3300.0,1638.1,494.36,3182.9,1686.6,0.0000,6725.6,4449.7,4252.8,3658.0,0.0000,-727.33,-262.02,-108.27,-72.187,-102.09,-587.69,0.0000,-1111.6,-1823.2,-743.89,-1533.5
152.0000000000,41687.,4669.1,8299.0,8155.7,4500.0,6017.1,13293.,1894.3,10542.,3086.1,5032.5,4280.7,0.0000,-11751.,-8690.2,-2078.2,-3813.3,-5204.1,-19414.,-371.68,-22288.,-6350.7,-4521.0,-3242.4,101.29,3608.3,3290.1,1635.2,492.91,3178.9,1686.6,0.0000,6723.3,4449.7,4252.8,3658.0,0.0000,-724.75,-260.90,-108.01,-71.952,-102.04,-587.69,0.0000,-1111.4,-1822.3,-744.12,-1532.7
153.0000000000,41592.,4622.6,8238.7,8156.0,4180.7,6019.9,13217.,1887.9,10481.,3086.9,5014.6,4242.3,0.0000,-11735.,-8685.8,-2078.2,-3809.0,-5198.0,-19403.,-370.67,-22279.,-6352.4,-4522.0,-3244.2,100.97,3597.0,3279.8,1632.3,491.41,3174.8,1686.6,0.0000,6720.8,4449.7,4252.8,3658.0,0.0000,-722.06,-259.76,-107.75,-71.707,-101.99,-587.69,0.0000,-1111.2,-1821.4,-744.35,-1532.0
154.0000000000,41494.,4494.7,8144.0,8103.8,3923.5,5972.4,13185.,1887.9,10427.,3057.5,4974.1,4229.2,0.0000,-11717.,-8681.1,-2078.1,-3804.6,-5191.9,-19393.,-369.70,-22270.,-6354.0,-4522.9,-3246.0,100.74,3588.8,3272.4,1631.1,490.34,3174.3,1686.6,0.0000,6720.6,4449.7,4252.8,3658.0,0.0000,-720.01,-258.83,-107.59,-71.525,-102.05,-587.69,0.0000,-1111.0,-1820.6,-744.58,-1531.2
155.0000000000,41493.,4389.0,8088.7,8002.8,3878.0,5878.5,13130.,1874.4,10387.,3024.7,4934.6,4185.7,0.0000,-11699.,-8676.3,-2077.9,-3800.3,-5185.7,-19382.,-368.73,-22261.,-6355.7,-4523.9,-3247.8,100.41,3577.2,3261.8,1628.1,488.79,3170.1,1686.6,0.0000,6718.1,4449.7,4252.8,3658.0,0.0000,-717.24,-257.65,-107.32,-71.273,-101.99,-587.69,0.0000,-1110.8,-1819.7,-744.79,-1530.4
156.0000000000,41435.,4382.4,8080.8,7948.7,3752.0,5877.4,13065.,1870.3,10343.,3022.3,4927.6,4159.0,0.0000,-11681.,-8671.3,-2077.7,-3795.9,-5179.5,-19371.,-367.76,-22252.,-6357.3,-4524.8,-3249.5,100.07,3564.9,3250.6,1624.8,487.15,3165.5,1686.6,0.0000,6715.4,4449.7,4252.8,3658.0,0.0000,-714.34,-256.42,-107.03,-71.007,-101.91,-587.69,0.0000,-1110.6,-1818.9,-745.00,-1529.6
157.0000000000,41175.,4341.9,8073.1,7890.0,3516.1,5882.8,12940.,1828.3,10307.,3020.6,4927.4,4153.0,0.0000,-11663.,-8666.2,-2077.4,-3791.5,-5173.2,-19360.,-366.80,-22243.,-6358.9,-4525.7,-3251.2,99.727,3552.7,3239.5,1621.5,485.52,3160.9,1686.6,0.0000,6712.7,4449.7,4252.8,3658.0,0.0000,-711.44,-255.18,-106.74,-70.743,-101.84,-587.69,0.0000,-1110.3,-1818.0,-745.21,-1528.8
158.0000000000,41080.,4300.5,6977.6,7838.5,3479.0,5797.3,12917.,1788.6,10306.,3021.4,4914.0,4139.4,0.0000,-11644.,-8660.8,-2077.0,-3787.1,-5166.8,-19349.,-365.85,-22234.,-6360.5,-4526.6,-3252.8,99.403,3541.2,3229.0,1618.5,483.98,3156.6,1686.6,0.0000,6710.1,4449.7,4252.8,3658.0,0.0000,-708.67,-253.99,-106.47,-70.491,-101.77,-587.69,0.0000,-1110.1,-1817.1,-745.41,-1528.0
159.0000000000,40950.,4298.0,6845.2,7742.6,3433.4,5676.8,12813.,1770.6,10306.,3011.8,4898.3,4118.1,0.0000,-11625.,-8655.5,-2076.6,-3782.7,-5160.4,-19339.,-365.08,-22225.,-6362.1,-4527.5,-3254.5,160.92,3564.1,3271.3,1623.2,492.24,3163.5,1686.6,0.0000,6714.2,4449.7,4252.8,3658.0,0.0000,-711.64,-255.43,-106.88,-70.853,-102.06,-587.69,0.0000,-1110.0,-1816.3,-745.61,-1527.3
160.0000000000,40837.,4300.0,6790.7,7667.7,3287.7,5561.6,12803.,1762.9,10305.,2968.8,4889.6,4095.9,0.0000,-11607.,-8650.5,-2076.3,-3778.4,-5154.0,-19328.,-364.10,-22217.,-6363.7,-4528.4,-3256.1,99.682,3551.1,3238.0,1620.9,485.30,3159.7,1686.6,0.0000,6711.9,4449.7,4252.8,3658.0,0.0000,-709.77,-254.00,-106.70,-70.649,-101.99,-587.69,0.0000,-1109.8,-1815.4,-745.81,-1526.5
161.0000000000,40749.,4240.6,6786.5,7668.3,3259.4,5480.0,12765.,1759.2,10185.,2954.5,4876.2,4083.5,0.0000,-11588.,-8645.4,-2075.9,-3774.1,-5147.6,-19317.,-363.11,-22208.,-6365.2,-4529.2,-3257.5,99.424,3541.9,3229.7,1618.1,484.07,3155.4,1686.6,0.0000,6709.4,4449.7,4252.8,3658.0,0.0000,-707.48,-252.99,-106.47,-70.447,-101.91,-587.69,0.0000,-1109.6,-1814.5,-746.01,-1525.7
162.0000000000,40681.,4194.8,6780.8,7667.9,3211.7,5461.6,12608.,1749.8,10165.,2935.4,4854.8,4084.4,0.0000,-11570.,-8640.1,-2075.5,-3769.7,-5141.2,-19307.,-362.14,-22199.,-6366.7,-4530.1,-3258.9,99.136,3531.7,3220.3,1615.1,482.70,3150.8,1686.6,0.0000,6706.6,4449.7,4252.8,3658.0,0.0000,-704.98,-251.89,-106.22,-70.222,-101.83,-587.69,0.0000,-1109.3,-1813.7,-746.20,-1524.9
163.0000000000,40637.,4064.7,6760.3,7543.1,3000.3,5459.3,12555.,1740.2,10131.,2936.2,4814.9,4081.3,0.0000,-11551.,-8634.6,-2075.1,-3765.4,-5134.8,-19296.,-361.18,-22190.,-6368.1,-4530.9,-3260.2,98.835,3520.9,3210.5,1612.0,481.26,3146.2,1686.6,0.0000,6703.9,4449.7,4252.8,3658.0,0.0000,-702.38,-250.77,-105.96,-69.988,-101.73,-587.69,0.0000,-1109.0,-1812.8,-746.40,-1524.0
164.0000000000,39921.,4030.0,6699.9,7459.3,2999.6,5456.5,12431.,1740.3,10061.,2937.1,4789.5,4054.8,0.0000,-11532.,-8628.9,-2074.6,-3761.0,-5128.2,-19286.,-360.24,-22182.,-6369.6,-4531.6,-3261.5,98.527,3510.0,3200.5,1608.9,479.80,3141.6,1686.6,0.0000,6701.2,4449.7,4252.8,3658.0,0.0000,-699.73,-249.62,-105.69,-69.749,-101.64,-587.69,0.0000,-1108.8,-1811.9,-746.59,-1523.2
165.0000000000,39581.,3923.1,6693.8,7458.2,2926.1,5454.0,12385.,1732.0,10025.,2937.9,4755.4,4023.5,0.0000,-11513.,-8623.2,-2074.1,-3756.7,-5121.6,-19276.,-359.42,-22173.,-6371.1,-4532.4,-3262.9,98.394,3505.2,3196.2,1609.2,479.19,3143.9,1686.6,1.5275,6702.9,4450.0,4252.8,3658.0,0.0000,-698.32,-248.91,-105.64,-69.634,-101.77,-587.69,-0.70100E-01,-1108.6,-1811.1,-746.77,-1522.4
166.0000000000,39454.,3910.3,6711.5,7458.2,2820.9,5455.9,12365.,1704.7,10004.,2938.8,4663.2,3969.1,0.0000,-11496.,-8618.5,-2073.8,-3752.6,-5115.1,-19265.,-359.55,-22165.,-6373.2,-4533.2,-3265.2,300.91,3715.9,3415.0,1656.7,505.87,3219.2,1686.6,70.321,6749.9,4456.4,4258.4,3664.2,0.0000,-721.69,-259.37,-108.75,-72.047,-104.15,-587.69,-3.2272,-1109.0,-1810.3,-746.99,-1522.2
167.0000000000,38931.,3907.5,6754.0,7465.5,2760.1,5465.5,12307.,1704.8,9941.1,2939.5,4611.3,3934.8,0.0000,-11484.,-8616.2,-2073.9,-3748.9,-5108.9,-19255.,-358.48,-22156.,-6374.8,-4533.9,-3266.5,102.72,3659.2,3336.6,1659.4,500.93,3222.6,1686.6,0.0000,6750.4,4451.1,4254.5,3659.1,0.0000,-728.24,-259.27,-109.51,-72.678,-104.42,-587.69,0.0000,-1108.9,-1809.4,-747.15,-1520.9
168.0000000000,38256.,3840.7,6722.3,7477.5,2694.3,5469.2,12146.,1695.2,9944.2,2940.1,4573.9,3915.0,0.0000,-11473.,-8614.2,-2074.0,-3745.2,-5103.0,-19245.,-357.24,-22148.,-6376.2,-4534.6,-3267.3,102.70,3658.6,3336.1,1657.0,500.29,3218.0,1686.6,0.0000,6747.2,4450.4,4253.6,3658.5,0.0000,-727.78,-258.97,-109.45,-72.651,-104.35,-587.69,0.0000,-1108.6,-1808.6,-747.33,-1520.1
169.0000000000,37403.,3836.8,6677.0,7473.1,2676.7,5411.8,12105.,1668.6,9944.1,2936.3,4547.4,3877.6,0.0000,-11462.,-8612.0,-2074.2,-3741.5,-5097.2,-19235.,-356.16,-22140.,-6377.5,-4535.4,-3268.1,102.73,3659.7,3337.0,1654.9,499.97,3213.3,1686.6,0.0000,6744.0,4449.8,4253.0,3658.1,0.0000,-727.67,-258.79,-109.42,-72.657,-104.34,-587.69,0.0000,-1108.4,-1807.7,-747.51,-1519.2
170.0000000000,36121.,3840.0,6637.4,7367.8,2676.9,5414.3,12043.,1668.7,9888.1,2937.2,4516.7,3844.7,0.0000,-11451.,-8609.3,-2074.3,-3737.8,-5091.2,-19225.,-355.12,-22131.,-6378.9,-4536.1,-3268.9,102.53,3652.7,3330.7,1652.2,498.94,3208.8,1686.6,0.0000,6741.2,4449.7,4252.8,3658.0,0.0000,-725.96,-258.04,-109.23,-72.505,-104.43,-587.69,0.0000,-1108.1,-1806.8,-747.69,-1518.4
171.0000000000,36072.,3837.9,6586.5,7354.4,2676.5,5415.2,12007.,1652.0,9853.0,2938.1,4493.3,3803.3,0.0000,-11439.,-8606.3,-2074.4,-3733.9,-5085.0,-19215.,-354.12,-22123.,-6380.3,-4536.8,-3269.7,102.22,3641.7,3320.6,1648.9,497.45,3203.9,1686.6,0.0000,6738.3,4449.7,4252.8,3658.0,0.0000,-723.43,-257.00,-108.96,-72.270,-104.49,-587.69,0.0000,-1107.9,-1806.0,-747.86,-1517.6
172.0000000000,35736.,3834.9,6523.3,7318.2,2675.6,5416.5,11981.,1632.7,9800.8,2939.0,4475.8,3802.0,0.0000,-11426.,-8602.9,-2074.4,-3730.0,-5078.7,-19205.,-353.17,-22115.,-6381.8,-4537.5,-3270.6,101.89,3629.8,3309.7,1645.5,495.86,3198.9,1686.6,0.0000,6735.3,4449.7,4252.8,3658.0,0.0000,-720.72,-255.89,-108.68,-72.017,-104.54,-587.69,0.0000,-1107.6,-1805.1,-748.04,-1516.7
173.0000000000,35694.,3789.7,6507.4,7218.6,2674.6,5407.3,11982.,1630.7,9749.4,2939.8,4459.3,3802.9,0.0000,-11412.,-8599.1,-2074.3,-3726.0,-5072.3,-19195.,-352.25,-22106.,-6383.2,-4538.1,-3271.4,101.54,3617.3,3298.4,1642.1,494.20,3193.8,1686.6,0.0000,6732.3,4449.7,4252.8,3658.0,0.0000,-717.90,-254.74,-108.38,-71.753,-104.59,-587.69,0.0000,-1107.4,-1804.2,-748.21,-1515.9
174.0000000000,35368.,3756.9,6499.0,7201.6,2620.3,5309.0,11911.,1606.3,9752.4,2936.7,4444.7,3803.7,0.0000,-11397.,-8594.9,-2074.0,-3722.0,-5065.8,-19186.,-351.37,-22098.,-6384.6,-4538.8,-3272.2,101.18,3604.6,3286.8,1638.5,492.49,3188.6,1686.6,0.0000,6729.2,4449.7,4252.8,3658.0,0.0000,-715.00,-253.56,-108.07,-71.482,-104.63,-587.69,0.0000,-1107.1,-1803.3,-748.38,-1515.1
175.0000000000,35210.,3746.0,6491.7,7079.4,2572.7,5277.3,11808.,1596.7,9740.8,2936.6,4440.2,3804.6,0.0000,-11382.,-8590.6,-2073.6,-3718.0,-5059.3,-19176.,-350.49,-22090.,-6386.0,-4539.5,-3273.0,100.82,3591.7,3275.0,1634.9,490.77,3183.4,1686.6,0.0000,6726.1,4449.7,4252.8,3658.0,0.0000,-712.05,-252.36,-107.76,-71.207,-104.66,-587.69,0.0000,-1106.9,-1802.4,-748.55,-1514.2
176.0000000000,34854.,3674.5,6483.2,7017.6,2536.7,5176.5,11766.,1583.6,9682.9,2928.9,4440.0,3789.9,0.0000,-11366.,-8586.0,-2073.1,-3713.9,-5052.6,-19166.,-349.63,-22081.,-6387.4,-4540.1,-3273.7,100.45,3578.6,3263.1,1631.3,489.02,3178.1,1686.6,0.0000,6723.0,4449.7,4252.8,3658.0,0.0000,-709.07,-251.14,-107.45,-70.929,-104.68,-587.69,0.0000,-1106.6,-1801.6,-748.72,-1513.4
177.0000000000,33940.,3609.0,6475.7,7015.9,2443.1,5112.2,11643.,1574.2,9655.6,2913.3,4428.9,3752.1,0.0000,-11350.,-8581.2,-2072.5,-3709.8,-5046.0,-19157.,-348.77,-22073.,-6388.8,-4540.8,-3274.4,100.08,3565.2,3250.9,1627.6,487.24,3172.6,1686.6,0.0000,6719.7,4449.7,4252.8,3658.0,0.0000,-706.02,-249.89,-107.13,-70.644,-104.69,-587.69,0.0000,-1106.4,-1800.7,-748.88,-1512.6
178.0000000000,33503.,3485.6,6465.9,6995.4,2395.3,5053.4,11528.,1560.9,9597.8,2914.1,4421.0,3700.8,0.0000,-11333.,-8576.3,-2071.9,-3705.7,-5039.3,-19147.,-347.91,-22064.,-6390.2,-4541.4,-3275.1,99.693,3551.5,3238.4,1623.6,485.40,3166.8,1686.6,0.0000,6716.3,4449.7,4252.8,3658.0,0.0000,-702.89,-248.61,-106.80,-70.352,-104.69,-587.69,0.0000,-1106.1,-1799.9,-749.05,-1511.8
179.0000000000,31990.,3430.7,6455.6,6942.3,2339.6,5049.5,11529.,1546.9,9468.5,2914.8,4420.8,3687.8,0.0000,-11315.,-8571.1,-2071.3,-3701.6,-5032.5,-19138.,-347.06,-22056.,-6391.5,-4542.0,-3275.7,99.315,3538.1,3226.1,1619.8,483.60,3161.1,1686.6,0.0000,6712.9,4449.7,4252.8,3658.0,0.0000,-699.81,-247.35,-106.47,-70.066,-104.69,-587.69,0.0000,-1105.9,-1799.0,-749.21,-1510.9
180.0000000000,31297.,3373.2,6445.1,6879.4,2282.1,5046.6,11530.,1536.7,9365.1,2910.8,4420.7,3674.8,0.0000,-11298.,-8565.7,-2070.5,-3697.5,-5025.7,-19128.,-346.21,-22048.,-6392.9,-4542.6,-3276.3,98.925,3524.2,3213.4,1615.8,481.74,3155.0,1686.6,0.0000,6709.3,4449.7,4252.8,3658.0,0.0000,-696.64,-246.04,-106.13,-69.770,-104.67,-587.69,0.0000,-1105.6,-1798.1,-749.37,-1510.1
181.0000000000,31153.,3366.0,6437.0,6710.7,2216.5,5044.0,11498.,1524.9,9330.8,2911.7,4420.4,3664.3,0.0000,-11280.,-8560.2,-2069.8,-3693.4,-5018.9,-19119.,-345.52,-22039.,-6394.3,-4543.2,-3277.1,98.948,3547.5,3253.8,1625.0,489.20,3174.8,1686.6,43.950,6721.1,4454.7,4254.9,3660.9,0.0000,-696.44,-246.61,-106.36,-69.818,-105.42,-587.69,-2.0166,-1105.5,-1797.3,-749.54,-1509.6
182.0000000000,30225.,3361.8,6431.8,6691.0,2100.2,5043.5,11405.,1513.2,9296.3,2912.6,4370.3,3634.2,0.0000,-11262.,-8554.8,-2069.2,-3689.3,-5012.2,-19110.,-344.65,-22031.,-6395.7,-4543.8,-3277.7,98.685,3515.6,3205.6,1619.6,480.70,3167.7,1686.6,0.0000,6717.0,4449.7,4252.8,3658.0,0.0000,-694.11,-244.78,-106.14,-69.560,-105.46,-587.69,0.0000,-1105.3,-1796.4,-749.69,-1508.5
183.0000000000,29314.,3356.4,6426.9,6569.9,2032.6,5043.0,11395.,1506.8,9259.7,2902.1,4326.4,3607.4,0.0000,-11244.,-8549.3,-2068.5,-3685.2,-5005.5,-19100.,-343.80,-22023.,-6397.0,-4544.4,-3278.1,98.559,3511.1,3201.5,1619.3,480.12,3168.4,1686.6,0.0000,6717.4,4449.7,4252.8,3658.0,0.0000,-692.81,-244.13,-106.07,-69.452,-105.77,-587.69,0.0000,-1105.1,-1795.5,-749.85,-1507.7
184.0000000000,27750.,3292.9,6422.8,6374.9,2023.2,5041.8,11222.,1506.8,9259.1,2894.4,4302.4,3547.5,0.0000,-11227.,-8543.8,-2067.8,-3681.1,-4998.9,-19091.,-342.93,-22015.,-6398.3,-4545.0,-3278.5,98.266,3500.7,3192.0,1616.5,478.73,3164.3,1686.6,0.0000,6715.0,4449.7,4252.8,3658.0,0.0000,-690.33,-243.06,-105.82,-69.226,-105.95,-587.69,0.0000,-1104.9,-1794.7,-750.01,-1506.9
185.0000000000,27472.,3277.6,6415.8,6301.6,1973.2,4984.9,11137.,1472.3,9149.6,2879.9,4242.7,3512.8,0.0000,-11209.,-8538.2,-2067.1,-3677.0,-4992.2,-19082.,-342.06,-22006.,-6399.5,-4545.6,-3278.9,97.961,3489.8,3182.1,1613.5,477.28,3160.0,1686.6,0.0000,6712.5,4449.7,4252.8,3658.0,0.0000,-687.76,-241.97,-105.56,-68.992,-106.11,-587.69,0.0000,-1104.7,-1793.8,-750.16,-1506.1
186.0000000000,27253.,3269.4,6409.2,6254.8,1903.9,4965.8,11081.,1459.0,9119.9,2871.3,4229.5,3469.5,0.0000,-11191.,-8532.4,-2066.4,-3673.0,-4985.5,-19073.,-341.21,-21998.,-6400.8,-4546.1,-3279.3,97.641,3478.4,3171.7,1610.3,475.75,3155.2,1686.6,0.0000,6709.6,4449.7,4252.8,3658.0,0.0000,-685.09,-240.83,-105.29,-68.747,-106.24,-587.69,0.0000,-1104.4,-1792.9,-750.31,-1505.3
187.0000000000,27011.,3261.4,6401.8,6161.5,1891.9,4963.1,10958.,1452.4,9062.5,2872.1,4206.5,3442.6,0.0000,-11173.,-8526.5,-2065.7,-3668.8,-4978.7,-19064.,-340.37,-21990.,-6402.1,-4546.7,-3279.6,97.315,3466.8,3161.1,1606.9,474.20,3150.2,1686.6,0.0000,6706.6,4449.7,4252.8,3658.0,0.0000,-682.37,-239.68,-105.00,-68.497,-106.37,-587.69,0.0000,-1104.2,-1792.1,-750.46,-1504.5
188.0000000000,26209.,3252.8,6392.6,6112.9,1881.7,4961.5,10934.,1452.5,9051.4,2855.6,4159.5,3416.2,0.0000,-11154.,-8520.5,-2064.9,-3664.7,-4971.9,-19055.,-339.53,-21982.,-6403.3,-4547.2,-3280.0,96.985,3455.1,3150.4,1603.5,472.63,3145.0,1686.6,0.0000,6703.5,4449.7,4252.8,3658.0,0.0000,-679.62,-238.51,-104.72,-68.245,-106.48,-587.69,0.0000,-1103.9,-1791.2,-750.61,-1503.7
189.0000000000,24998.,3244.4,6383.3,6020.7,1798.5,4959.4,10837.,1452.5,8970.2,2853.9,4141.2,3402.8,0.0000,-11136.,-8514.4,-2064.0,-3660.6,-4965.0,-19046.,-338.70,-21973.,-6404.6,-4547.8,-3280.4,96.652,3443.2,3139.6,1600.0,471.04,3139.6,1686.6,0.0000,6700.3,4449.7,4252.8,3658.0,0.0000,-676.85,-237.34,-104.43,-67.990,-106.57,-587.69,0.0000,-1103.7,-1790.3,-750.76,-1502.9
190.0000000000,23031.,3182.3,5998.1,5992.8,1760.6,4956.5,10664.,1452.5,8913.8,2854.8,4124.4,3386.7,0.0000,-11117.,-8508.2,-2063.1,-3656.5,-4958.0,-19037.,-337.88,-21965.,-6405.8,-4548.3,-3281.8,96.326,3431.6,3129.0,1596.5,469.48,3134.4,1686.6,0.0000,6697.2,4449.7,4252.8,3658.0,0.0000,-674.12,-236.18,-104.14,-67.741,-106.67,-587.69,0.0000,-1103.5,-1789.5,-750.91,-1502.2
191.0000000000,22780.,3144.7,5240.0,5922.8,1727.9,4953.0,10627.,1439.1,8912.4,2855.6,4102.6,3363.9,0.0000,-11098.,-8501.9,-2062.2,-3652.3,-4951.0,-19028.,-337.05,-21957.,-6407.0,-4548.8,-3283.5,95.998,3419.9,3118.4,1593.0,467.92,3129.0,1686.6,0.0000,6694.0,4449.7,4252.8,3658.0,0.0000,-671.38,-235.02,-103.85,-67.490,-106.75,-587.69,0.0000,-1103.2,-1788.6,-751.06,-1501.4
192.0000000000,22707.,3135.9,5231.1,5808.4,1694.5,4948.8,10577.,1416.2,8910.9,2856.4,4070.6,3354.3,0.0000,-11079.,-8495.5,-2061.2,-3648.2,-4944.0,-19020.,-336.23,-21949.,-6408.2,-4549.3,-3284.8,95.667,3408.1,3107.6,1589.4,466.33,3123.4,1686.6,0.0000,6690.7,4449.7,4252.8,3658.0,0.0000,-668.61,-233.84,-103.56,-67.237,-106.82,-587.69,0.0000,-1103.0,-1787.8,-751.20,-1500.6
193.0000000000,22409.,3196.2,5221.6,5668.2,1693.3,4944.4,10496.,1413.4,8908.9,2857.3,4061.2,3347.3,0.0000,-11060.,-8489.1,-2060.2,-3644.0,-4937.0,-19011.,-335.42,-21941.,-6409.4,-4549.8,-3285.7,95.335,3396.3,3096.8,1585.8,464.75,3117.8,1686.6,0.0000,6687.3,4449.7,4252.8,3658.0,0.0000,-665.85,-232.67,-103.27,-66.984,-106.89,-587.69,0.0000,-1102.8,-1786.9,-751.34,-1499.8
194.0000000000,22124.,3187.6,5212.2,5561.4,1683.0,4940.2,10408.,1380.0,8906.7,2858.1,4031.1,3348.2,0.0000,-11040.,-8482.6,-2059.1,-3639.9,-4929.9,-19002.,-334.60,-21932.,-6410.6,-4550.3,-3286.5,95.008,3384.6,3086.2,1582.3,463.19,3112.2,1686.6,0.0000,6684.0,4449.7,4252.8,3658.0,0.0000,-663.10,-231.50,-102.97,-66.733,-106.94,-587.69,0.0000,-1102.5,-1786.0,-751.49,-1499.0
195.0000000000,20447.,3178.8,5202.8,5460.2,1622.0,4945.1,10360.,1380.0,8882.0,2859.0,4026.2,3341.7,0.0000,-11021.,-8476.1,-2058.1,-3635.8,-4922.8,-18994.,-333.79,-21924.,-6411.7,-4550.8,-3287.2,94.689,3373.2,3075.8,1578.8,461.66,3106.7,1686.6,0.0000,6680.7,4449.7,4252.8,3658.0,0.0000,-660.42,-230.35,-102.69,-66.489,-107.00,-587.69,0.0000,-1102.3,-1785.2,-751.63,-1498.2
196.0000000000,19702.,3170.9,5194.1,5457.5,1562.6,4941.1,10326.,1376.5,8742.2,2859.8,3996.1,3309.6,0.0000,-11002.,-8469.6,-2057.0,-3631.6,-4915.7,-18985.,-333.02,-21916.,-6412.9,-4551.3,-3287.9,94.480,3365.8,3069.0,1577.1,460.67,3104.7,1686.6,0.0000,6679.5,4449.7,4252.8,3658.0,0.0000,-658.50,-229.48,-102.53,-66.322,-107.17,-587.69,0.0000,-1102.1,-1784.3,-751.77,-1497.4
197.0000000000,19696.,3179.4,5200.8,5455.5,1511.9,4939.0,10280.,1361.9,8624.5,2860.7,3972.9,3279.0,0.0000,-10984.,-8463.8,-2056.0,-3627.7,-4908.6,-18976.,-332.59,-21908.,-6414.3,-4551.8,-3289.0,126.65,3465.4,3167.8,1603.5,475.32,3145.9,1686.6,24.827,6704.7,4453.4,4255.2,3660.7,0.0000,-672.57,-234.84,-104.40,-67.794,-108.77,-587.69,-1.1389,-1102.2,-1783.5,-751.92,-1496.9
198.0000000000,19697.,3209.3,5227.9,5390.1,1440.9,4942.1,10104.,1361.9,8623.7,2861.5,3971.8,3267.6,0.0000,-10970.,-8459.8,-2055.3,-3624.0,-4901.7,-18968.,-331.92,-21900.,-6415.6,-4552.3,-3289.9,272.84,3615.5,3342.8,1630.9,496.87,3182.2,1686.6,107.59,6731.4,4466.3,4267.4,3672.5,0.0000,-680.02,-240.17,-105.40,-68.662,-109.88,-587.69,-4.9356,-1102.2,-1782.7,-752.11,-1497.3
199.0000000000,18785.,3233.4,5251.5,5333.8,1445.7,4948.7,9928.7,1362.0,8524.1,2835.7,3970.7,3229.4,0.0000,-10957.,-8456.6,-2054.8,-3620.5,-4895.0,-18960.,-331.03,-21892.,-6416.7,-4552.7,-3290.2,98.263,3500.6,3191.9,1617.7,478.74,3167.4,1686.6,0.0000,6716.9,4449.7,4252.8,3658.0,0.0000,-683.69,-237.75,-105.86,-68.940,-110.10,-587.69,0.0000,-1102.0,-1781.8,-752.18,-1495.2
200.0000000000,17942.,3250.2,5268.8,5204.4,1449.0,4954.6,9872.9,1362.0,8291.4,2823.7,3947.0,3222.3,0.0000,-10946.,-8453.7,-2054.4,-3617.0,-4888.6,-18951.,-330.16,-21884.,-6417.7,-4553.2,-3290.5,136.97,3603.2,3326.9,1620.3,480.64,3169.7,1686.6,0.0000,6718.2,4449.7,4252.8,3658.0,0.0000,-686.38,-241.07,-106.16,-69.214,-110.42,-587.69,0.0000,-1101.9,-1781.0,-752.32,-1494.5
201.0000000000,17554.,3260.5,5279.3,5188.4,1450.6,4954.9,9785.1,1362.0,8282.2,2814.8,3934.3,3190.8,0.0000,-10935.,-8450.9,-2054.1,-3613.6,-4882.2,-18943.,-329.26,-21876.,-6418.8,-4553.6,-3290.7,98.683,3515.5,3205.6,1618.7,480.68,3165.4,1686.6,0.0000,6715.6,4449.7,4252.8,3658.0,0.0000,-685.95,-238.26,-106.11,-69.214,-110.50,-587.69,0.0000,-1101.7,-1780.2,-752.45,-1493.7
202.0000000000,17413.,3264.0,5284.9,5021.0,1420.5,4888.2,9601.4,1362.1,8257.5,2796.6,3926.4,3173.9,0.0000,-10924.,-8448.0,-2053.7,-3610.1,-4875.6,-18934.,-328.41,-21869.,-6419.8,-4554.1,-3291.0,98.630,3513.6,3203.9,1616.9,480.41,3161.3,1686.6,0.0000,6713.1,4449.7,4252.8,3658.0,0.0000,-685.26,-237.89,-106.02,-69.165,-110.58,-587.69,0.0000,-1101.4,-1779.3,-752.57,-1493.0
203.0000000000,17392.,3265.3,5287.8,4935.3,1387.2,4888.5,9446.9,1362.0,8185.2,2786.6,3886.2,3165.6,0.0000,-10914.,-8444.8,-2053.2,-3606.5,-4869.0,-18926.,-327.59,-21861.,-6420.8,-4554.6,-3291.2,98.425,3506.3,3197.2,1614.4,479.42,3157.1,1686.6,0.0000,6710.6,4449.7,4252.8,3658.0,0.0000,-683.51,-237.14,-105.83,-69.007,-110.66,-587.69,0.0000,-1101.2,-1778.5,-752.67,-1492.2
204.0000000000,17337.,3262.9,5285.8,4936.1,1355.7,4890.1,9278.7,1362.0,8185.8,2787.5,3878.4,3118.2,0.0000,-10902.,-8441.4,-2052.7,-3602.9,-4862.2,-18918.,-326.77,-21853.,-6421.8,-4555.2,-3291.4,98.154,3496.7,3188.4,1611.3,478.13,3152.1,1686.6,0.0000,6707.6,4449.7,4252.8,3658.0,0.0000,-681.31,-236.24,-105.59,-68.804,-110.70,-587.69,0.0000,-1101.0,-1777.6,-752.77,-1491.4
205.0000000000,17061.,3258.9,5263.2,4935.5,1322.0,4892.4,9150.7,1362.1,8190.4,2788.3,3878.3,3096.8,0.0000,-10891.,-8437.6,-2052.1,-3599.3,-4855.3,-18910.,-325.97,-21846.,-6422.8,-4555.9,-3291.7,97.859,3486.2,3178.8,1608.0,476.72,3147.0,1686.6,0.0000,6704.6,4449.7,4252.8,3658.0,0.0000,-678.93,-235.27,-105.32,-68.582,-110.73,-587.69,0.0000,-1100.8,-1776.7,-752.86,-1490.7
206.0000000000,16316.,3254.0,5205.8,4881.9,1320.9,4900.2,9057.7,1360.1,8192.2,2781.4,3844.1,3086.4,0.0000,-10879.,-8433.7,-2051.3,-3595.6,-4848.4,-18902.,-325.18,-21838.,-6423.8,-4556.7,-3291.9,97.544,3475.0,3168.6,1604.6,475.21,3141.6,1686.6,0.0000,6701.4,4449.7,4252.8,3658.0,0.0000,-676.40,-234.25,-105.04,-68.345,-110.76,-587.69,0.0000,-1100.6,-1775.9,-752.95,-1489.9
207.0000000000,16236.,3231.0,5198.9,4728.9,1319.7,4900.4,8984.6,1343.9,8139.4,2765.0,3821.8,3087.2,0.0000,-10866.,-8429.5,-2050.5,-3592.0,-4841.5,-18894.,-324.40,-21830.,-6424.8,-4557.5,-3292.1,97.219,3463.4,3158.0,1601.1,473.66,3136.1,1686.6,0.0000,6698.1,4449.7,4252.8,3658.0,0.0000,-673.78,-233.20,-104.76,-68.101,-110.77,-587.69,0.0000,-1100.4,-1775.0,-753.05,-1489.2
208.0000000000,16158.,3224.8,5192.9,4726.7,1228.7,4897.4,8775.6,1344.0,8122.3,2765.9,3813.8,3087.9,0.0000,-10854.,-8425.2,-2049.6,-3588.3,-4834.5,-18885.,-323.64,-21822.,-6425.8,-4558.2,-3292.3,96.999,3455.6,3150.9,1598.8,472.61,3132.6,1686.6,0.0000,6696.0,4449.7,4252.8,3658.0,0.0000,-671.90,-232.39,-104.56,-67.930,-110.85,-587.69,0.0000,-1100.2,-1774.2,-753.14,-1488.4
209.0000000000,16117.,3287.8,5186.5,4635.4,1189.7,4893.7,8716.6,1339.6,8088.8,2766.7,3796.7,3071.9,0.0000,-10841.,-8420.8,-2048.7,-3584.6,-4827.5,-18877.,-322.87,-21815.,-6426.8,-4558.9,-3292.5,96.677,3444.1,3140.4,1595.3,471.07,3127.3,1686.6,0.0000,6692.9,4449.7,4252.8,3658.0,0.0000,-669.29,-231.34,-104.28,-67.687,-110.85,-587.69,0.0000,-1099.9,-1773.3,-753.23,-1487.6
210.0000000000,16047.,3280.9,5178.4,4586.0,1188.6,4889.9,8538.2,1319.5,8009.1,2767.6,3784.5,3062.5,0.0000,-10828.,-8416.3,-2047.7,-3580.9,-4820.5,-18869.,-322.15,-21807.,-6427.7,-4559.5,-3292.7,96.390,3433.9,3131.1,1594.3,469.74,3129.8,1686.6,4.0811,6695.8,4451.0,4255.6,3658.2,0.0000,-666.90,-230.40,-104.10,-67.470,-111.09,-587.69,-0.18718,-1099.8,-1772.5,-753.34,-1486.9
211.0000000000,15994.,3269.4,5170.2,4580.7,1187.4,4887.2,8449.5,1307.9,7925.1,2768.4,3784.4,3028.8,0.0000,-10815.,-8411.6,-2046.8,-3577.1,-4813.6,-18862.,-321.39,-21799.,-6428.7,-4560.2,-3292.9,96.053,3421.8,3120.1,1590.7,468.13,3122.2,1686.6,0.0000,6689.9,4449.7,4252.8,3658.0,0.0000,-664.14,-229.34,-103.80,-67.216,-111.06,-587.69,0.0000,-1099.6,-1771.6,-753.42,-1486.1
212.0000000000,15972.,3248.6,5161.1,4453.4,1186.1,4804.1,8325.7,1307.9,7893.4,2769.3,3784.4,3010.8,0.0000,-10801.,-8406.7,-2045.7,-3573.4,-4806.6,-18854.,-320.64,-21791.,-6429.6,-4560.8,-3293.0,95.714,3409.7,3109.1,1587.0,466.51,3116.5,1686.6,0.0000,6686.5,4449.7,4252.8,3658.0,0.0000,-661.36,-228.27,-103.50,-66.961,-111.04,-587.69,0.0000,-1099.3,-1770.8,-753.51,-1485.4
213.0000000000,15656.,3240.2,5151.6,4444.6,1184.8,4738.6,8299.0,1307.8,7891.3,2770.1,3784.3,2976.9,0.0000,-10787.,-8401.6,-2044.7,-3569.6,-4799.6,-18846.,-319.90,-21784.,-6430.5,-4561.4,-3293.1,95.370,3397.5,3097.9,1583.2,464.86,3110.5,1686.6,0.0000,6682.9,4449.7,4252.8,3658.0,0.0000,-658.54,-227.18,-103.19,-66.702,-111.00,-587.69,0.0000,-1099.1,-1770.0,-753.59,-1484.6
214.0000000000,14603.,3231.4,5142.4,4390.7,1178.9,4734.8,8254.4,1274.3,7831.0,2770.8,3784.2,2949.1,0.0000,-10773.,-8396.4,-2043.6,-3565.9,-4792.6,-18838.,-319.17,-21776.,-6431.4,-4562.0,-3293.2,95.024,3385.2,3086.7,1579.3,463.21,3104.4,1686.6,0.0000,6679.2,4449.7,4252.8,3658.0,0.0000,-655.71,-226.09,-102.88,-66.443,-110.96,-587.69,0.0000,-1098.9,-1769.1,-753.68,-1483.9
215.0000000000,14269.,3176.8,5134.0,4340.3,1117.8,4714.8,8190.9,1234.2,7784.2,2752.0,3784.0,2948.8,0.0000,-10759.,-8391.0,-2042.4,-3562.1,-4785.5,-18830.,-318.45,-21768.,-6432.2,-4562.5,-3293.2,94.677,3372.8,3075.5,1575.4,461.55,3098.2,1686.6,0.0000,6675.5,4449.7,4252.8,3658.0,0.0000,-652.85,-224.98,-102.57,-66.182,-110.91,-587.69,0.0000,-1098.7,-1768.3,-753.77,-1483.1
216.0000000000,14233.,3148.6,5125.5,4270.8,1116.5,4644.2,8075.7,1218.0,7747.7,2752.8,3777.1,2946.4,0.0000,-10744.,-8385.5,-2041.3,-3558.3,-4778.4,-18822.,-317.75,-21760.,-6433.1,-4563.1,-3293.2,94.336,3360.7,3064.4,1571.6,459.92,3092.1,1686.6,0.0000,6671.9,4449.7,4252.8,3658.0,0.0000,-650.03,-223.89,-102.26,-65.925,-110.85,-587.69,0.0000,-1098.5,-1767.5,-753.86,-1482.4
217.0000000000,13311.,3139.7,5116.0,4200.7,1115.2,4632.7,7934.6,1200.0,7746.0,2753.6,3741.5,2904.4,0.0000,-10729.,-8379.9,-2040.0,-3554.5,-4771.3,-18815.,-317.04,-21753.,-6434.0,-4563.6,-3293.2,93.997,3348.6,3053.4,1567.8,458.30,3085.9,1686.6,0.0000,6668.2,4449.7,4252.8,3658.0,0.0000,-647.22,-222.80,-101.96,-65.670,-110.79,-587.69,0.0000,-1098.3,-1766.7,-753.95,-1481.6
218.0000000000,13067.,3130.7,4139.2,4159.5,1113.8,4628.3,7642.0,1187.9,7744.0,2754.4,3713.0,2896.8,0.0000,-10714.,-8374.1,-2038.8,-3550.7,-4764.2,-18807.,-316.34,-21745.,-6434.8,-4564.2,-3293.2,93.660,3336.6,3042.4,1563.9,456.69,3079.7,1686.6,0.0000,6664.5,4449.7,4252.8,3658.0,0.0000,-644.42,-221.71,-101.66,-65.416,-110.73,-587.69,0.0000,-1098.1,-1765.9,-754.03,-1480.9
219.0000000000,12985.,3121.7,3974.7,4147.5,1112.5,4623.9,7589.4,1182.0,7724.9,2755.2,3690.9,2882.2,0.0000,-10699.,-8368.2,-2037.5,-3546.9,-4757.1,-18799.,-315.65,-21737.,-6435.6,-4564.7,-3293.2,93.324,3324.6,3031.5,1560.1,455.08,3073.5,1686.6,0.0000,6660.8,4449.7,4252.8,3658.0,0.0000,-641.62,-220.62,-101.35,-65.163,-110.65,-587.69,0.0000,-1097.9,-1765.1,-754.12,-1480.2
220.0000000000,11918.,3112.7,3965.5,3960.6,1101.8,4619.3,7493.2,1182.0,7601.8,2756.0,3672.3,2860.4,0.0000,-10684.,-8362.2,-2036.2,-3543.1,-4749.9,-18792.,-314.95,-21729.,-6436.5,-4565.2,-3293.1,92.988,3312.7,3020.6,1556.2,453.47,3067.2,1686.6,0.0000,6657.1,4449.7,4252.8,3658.0,0.0000,-638.82,-219.53,-101.05,-64.910,-110.57,-587.69,0.0000,-1097.7,-1764.3,-754.20,-1479.4
221.0000000000,11525.,3103.7,3956.0,3944.1,1045.8,4614.1,7441.6,1182.0,7599.7,2756.8,3636.8,2831.0,0.0000,-10668.,-8356.2,-2034.8,-3539.3,-4742.7,-18784.,-314.25,-21722.,-6437.3,-4565.7,-3293.0,92.656,3300.8,3009.8,1552.3,451.88,3061.0,1686.6,0.0000,6653.3,4449.7,4252.8,3658.0,0.0000,-636.05,-218.45,-100.74,-64.660,-110.49,-587.69,0.0000,-1097.5,-1763.5,-754.29,-1478.7
222.0000000000,11525.,3094.8,3946.5,3940.8,1044.5,4609.0,7394.0,1182.1,7504.2,2757.5,3635.1,2810.6,0.0000,-10652.,-8350.1,-2033.5,-3535.5,-4735.5,-18777.,-313.56,-21714.,-6438.1,-4566.2,-3292.9,92.337,3289.4,2999.4,1548.6,450.35,3054.9,1686.6,0.0000,6649.7,4449.7,4252.8,3658.0,0.0000,-633.35,-217.40,-100.45,-64.419,-110.41,-587.69,0.0000,-1097.2,-1762.7,-754.37,-1478.0
223.0000000000,11476.,3035.9,3937.2,3937.3,1043.3,4603.8,7335.9,1182.1,7457.7,2758.3,3635.0,2780.2,0.0000,-10637.,-8344.0,-2032.1,-3531.7,-4728.2,-18769.,-312.87,-21706.,-6438.9,-4566.7,-3292.8,92.036,3278.7,2989.6,1545.1,448.91,3049.1,1686.6,0.0000,6646.2,4449.7,4252.8,3658.0,0.0000,-630.78,-216.38,-100.17,-64.190,-110.33,-587.69,0.0000,-1097.0,-1761.9,-754.45,-1477.2
224.0000000000,10145.,3012.6,3928.3,3934.2,987.76,4598.6,7274.3,1166.1,7455.1,2759.1,3635.0,2750.3,0.0000,-10621.,-8337.8,-2030.6,-3527.9,-4720.9,-18762.,-312.20,-21699.,-6439.7,-4567.2,-3292.7,91.759,3268.9,2980.7,1542.5,447.60,3045.6,1686.6,0.0000,6644.2,4449.7,4252.8,3658.0,0.0000,-628.38,-215.43,-99.946,-63.979,-110.34,-587.69,0.0000,-1096.9,-1761.1,-754.54,-1476.5
225.0000000000,10061.,3004.7,3919.7,3843.9,914.06,4593.9,7218.9,1145.6,7452.4,2757.3,3634.9,2739.2,0.0000,-10605.,-8331.6,-2029.2,-3524.1,-4713.7,-18755.,-311.51,-21691.,-6440.4,-4567.6,-3292.6,91.459,3258.2,2970.9,1539.0,446.16,3039.8,1686.6,0.0000,6640.7,4449.7,4252.8,3658.0,0.0000,-625.81,-214.42,-99.671,-63.752,-110.26,-587.69,0.0000,-1096.7,-1760.4,-754.62,-1475.8
226.0000000000,8587.3,2968.5,3910.9,3754.1,912.82,4581.4,7082.2,1128.1,7397.3,2738.3,3624.5,2723.0,0.0000,-10588.,-8325.4,-2027.8,-3520.3,-4706.5,-18747.,-310.82,-21683.,-6441.2,-4568.1,-3292.4,91.154,3247.3,2961.0,1535.4,444.69,3033.9,1686.6,0.0000,6637.2,4449.7,4252.8,3658.0,0.0000,-623.21,-213.40,-99.390,-63.521,-110.16,-587.69,0.0000,-1096.5,-1759.6,-754.70,-1475.0
227.0000000000,8275.9,2919.3,3902.1,3653.6,911.60,4513.7,7022.0,1102.0,7367.4,2736.6,3601.7,2716.0,0.0000,-10572.,-8319.2,-2026.3,-3516.5,-4699.2,-18740.,-310.13,-21675.,-6442.0,-4568.6,-3292.3,90.853,3236.6,2951.2,1531.8,443.26,3028.0,1686.6,0.0000,6633.6,4449.7,4252.8,3658.0,0.0000,-620.65,-212.39,-99.114,-63.294,-110.07,-587.69,0.0000,-1096.3,-1758.8,-754.78,-1474.3
228.0000000000,8046.1,2911.1,3893.2,3650.6,871.10,4508.7,7005.5,1092.1,7306.2,2737.4,3597.8,2705.4,0.0000,-10556.,-8313.0,-2024.8,-3512.7,-4691.9,-18732.,-309.45,-21668.,-6442.7,-4569.0,-3292.1,90.559,3226.1,2941.7,1528.3,441.85,3022.1,1686.6,0.0000,6630.1,4449.7,4252.8,3658.0,0.0000,-618.12,-211.39,-98.842,-63.072,-109.97,-587.69,0.0000,-1096.1,-1758.1,-754.86,-1473.6
229.0000000000,7660.2,2903.1,3884.3,3642.5,845.21,4437.2,6939.5,1092.1,7303.2,2720.4,3592.6,2706.1,0.0000,-10539.,-8306.6,-2023.3,-3508.9,-4684.6,-18725.,-308.77,-21660.,-6443.4,-4569.4,-3291.9,90.273,3215.9,2932.4,1524.9,440.47,3016.5,1686.6,0.0000,6626.8,4449.7,4252.8,3658.0,0.0000,-615.65,-210.42,-98.578,-62.854,-109.88,-587.69,0.0000,-1096.1,-1757.3,-754.94,-1472.9
230.0000000000,7610.5,2895.4,3876.1,3536.2,844.05,4387.0,6840.4,1079.5,7296.7,2719.2,3579.1,2689.7,0.0000,-10523.,-8300.3,-2021.8,-3505.1,-4677.2,-18718.,-308.09,-21652.,-6444.2,-4569.9,-3291.7,89.989,3205.8,2923.2,1521.5,439.11,3010.8,1686.6,0.0000,6623.4,4449.7,4252.8,3658.0,0.0000,-613.20,-209.45,-98.315,-62.639,-109.78,-587.69,0.0000,-1096.0,-1756.6,-755.02,-1472.1
231.0000000000,7601.3,2887.9,3867.3,3437.1,842.94,4350.9,6816.3,1074.2,7293.3,2714.8,3569.8,2654.2,0.0000,-10506.,-8294.0,-2020.3,-3501.4,-4669.9,-18711.,-307.41,-21644.,-6444.9,-4570.3,-3291.5,89.712,3195.9,2914.2,1518.1,437.78,3005.2,1686.6,0.0000,6620.0,4449.7,4252.8,3658.0,0.0000,-610.79,-208.49,-98.058,-62.429,-109.68,-587.69,0.0000,-1095.9,-1755.8,-755.10,-1471.4
232.0000000000,7519.7,2880.8,3859.1,3434.0,791.59,4305.3,6733.4,1071.1,7282.3,2710.9,3551.0,2644.8,0.0000,-10490.,-8287.7,-2018.7,-3497.6,-4662.5,-18703.,-306.74,-21637.,-6445.6,-4570.7,-3291.2,89.438,3186.2,2905.3,1514.8,436.47,2999.7,1686.6,0.0000,6616.7,4449.7,4252.8,3658.0,0.0000,-608.41,-207.55,-97.803,-62.220,-109.57,-587.69,0.0000,-1095.8,-1755.0,-755.18,-1470.7
233.0000000000,7482.4,2873.6,3850.9,3431.0,776.62,4270.2,6571.4,1029.6,7219.6,2711.7,3541.7,2634.0,0.0000,-10473.,-8281.4,-2017.2,-3493.8,-4655.1,-18696.,-306.06,-21629.,-6446.3,-4571.1,-3291.0,89.168,3176.6,2896.5,1511.5,435.17,2994.2,1686.6,0.0000,6613.4,4449.7,4252.8,3658.0,0.0000,-606.05,-206.61,-97.552,-62.015,-109.47,-587.69,0.0000,-1095.8,-1754.3,-755.26,-1469.9
234.0000000000,7446.9,2866.3,3842.9,3428.0,775.54,4265.4,6499.6,1007.7,7216.8,2712.4,3541.6,2599.8,0.0000,-10457.,-8275.2,-2015.6,-3490.1,-4647.7,-18689.,-305.40,-21622.,-6447.0,-4571.5,-3290.7,88.904,3167.2,2887.9,1508.4,433.91,2989.2,1686.6,0.0000,6610.4,4449.7,4252.8,3658.0,0.0000,-603.74,-205.70,-97.312,-61.814,-109.38,-587.69,0.0000,-1095.7,-1753.5,-755.33,-1469.2
235.0000000000,7358.1,2859.2,3834.9,3384.0,728.08,4211.5,6443.5,1002.3,7098.5,2701.0,3541.5,2574.8,0.0000,-10440.,-8268.9,-2014.0,-3486.3,-4640.3,-18682.,-304.73,-21614.,-6447.7,-4571.9,-3290.4,88.645,3157.9,2879.5,1505.2,432.66,2983.9,1686.6,0.0000,6607.3,4449.7,4252.8,3658.0,0.0000,-601.46,-204.79,-97.070,-61.616,-109.28,-587.69,0.0000,-1095.6,-1752.8,-755.41,-1468.5
236.0000000000,7323.2,2859.9,3834.4,3286.4,710.62,4175.4,6287.0,1002.4,7055.6,2684.0,3541.4,2559.3,0.0000,-10424.,-8263.1,-2012.5,-3482.7,-4632.9,-18675.,-304.24,-21606.,-6448.5,-4572.3,-3290.4,95.937,3196.6,2913.3,1517.4,437.62,3002.7,1686.6,3.2382,6619.1,4451.0,4254.2,3659.2,0.0000,-607.71,-206.83,-97.957,-62.294,-110.03,-587.69,-0.14847,-1095.7,-1752.1,-755.49,-1467.9
237.0000000000,7005.0,2870.2,3842.6,3249.2,622.26,4112.4,6095.3,983.10,7053.6,2670.2,3529.3,2540.2,0.0000,-10410.,-8258.0,-2011.1,-3479.1,-4625.6,-18668.,-303.56,-21599.,-6449.2,-4572.7,-3290.1,89.715,3196.1,2914.3,1516.3,437.77,3000.6,1686.6,0.0000,6617.2,4449.7,4252.9,3658.0,0.0000,-607.74,-206.69,-97.999,-62.332,-110.08,-587.69,0.0000,-1095.7,-1751.4,-755.56,-1467.0
238.0000000000,6909.5,2873.9,3846.1,3218.8,584.80,4111.8,5798.7,966.54,7048.7,2669.9,3522.7,2520.9,0.0000,-10396.,-8253.2,-2009.8,-3475.7,-4618.4,-18661.,-302.88,-21591.,-6449.9,-4573.0,-3289.7,89.710,3195.9,2914.1,1515.9,437.74,2999.6,1686.6,0.0000,6616.6,4449.7,4252.8,3660.6,0.0000,-607.23,-206.40,-97.983,-62.315,-110.13,-587.69,0.0000,-1095.6,-1750.7,-755.64,-1466.6
239.0000000000,6849.8,2887.8,3859.1,3219.5,524.18,4112.6,5570.5,953.85,7034.1,2666.7,3522.6,2476.2,0.0000,-10383.,-8249.0,-2008.6,-3472.3,-4611.3,-18654.,-302.41,-21584.,-6450.7,-4573.4,-3289.6,191.32,3339.6,3000.7,1555.0,449.75,3060.7,1686.6,64.743,6657.8,4462.3,4265.6,3674.0,0.0000,-620.89,-211.32,-100.01,-63.751,-112.17,-587.69,-2.9683,-1096.0,-1750.0,-755.77,-1467.0
240.0000000000,6847.6,2882.1,3893.9,3225.3,529.66,4120.1,5467.8,908.84,7028.3,2667.4,3520.4,2459.2,0.0000,-10374.,-8246.6,-2007.8,-3469.3,-4604.5,-18647.,-301.88,-21577.,-6451.5,-4573.8,-3289.5,336.87,3824.5,3421.4,1614.5,472.78,3149.3,1686.6,324.54,6724.6,4486.7,4292.3,3703.2,0.0000,-634.37,-223.17,-102.11,-65.171,-114.85,-587.69,-14.879,-1096.5,-1749.3,-755.96,-1468.9
241.0000000000,6811.3,2894.7,3929.7,3237.8,535.83,4135.1,5403.1,894.55,7004.9,2668.0,3497.8,2417.0,0.0000,-10367.,-8245.5,-2007.4,-3466.5,-4598.1,-18640.,-301.14,-21570.,-6452.1,-4574.1,-3289.0,94.435,3364.2,3067.6,1599.3,468.86,3130.0,1686.6,0.0000,6708.2,4455.0,4261.7,3660.3,0.0000,-638.03,-216.65,-102.69,-65.636,-114.98,-587.69,0.0000,-1096.4,-1748.6,-755.90,-1464.5
242.0000000000,6786.0,2914.7,3952.0,3203.0,539.90,4148.9,5187.6,876.68,6947.7,2668.8,3485.5,2403.1,0.0000,-10361.,-8244.6,-2007.1,-3463.8,-4592.2,-18633.,-300.39,-21563.,-6452.6,-4574.5,-3288.5,94.453,3364.8,3068.2,1584.5,462.59,3120.1,1686.6,0.0000,6690.7,4450.3,4253.7,3658.1,0.0000,-637.82,-216.53,-102.70,-65.599,-115.01,-587.69,0.0000,-1096.3,-1748.0,-755.94,-1463.6
243.0000000000,6723.3,2922.1,3960.9,3145.1,541.05,4093.4,5151.6,876.70,6943.5,2669.4,3485.4,2379.8,0.0000,-10354.,-8243.2,-2006.9,-3460.9,-4586.3,-18626.,-299.67,-21556.,-6453.1,-4574.8,-3287.9,94.324,3360.2,3064.0,1581.9,460.57,3118.0,1686.6,0.0000,6688.1,4449.7,4252.9,3658.0,0.0000,-636.63,-216.07,-102.60,-65.492,-115.06,-587.69,0.0000,-1096.2,-1747.3,-756.01,-1462.9
244.0000000000,6466.0,2923.2,3962.9,3061.5,540.73,4094.7,5102.8,873.53,6946.4,2670.1,3478.2,2365.4,0.0000,-10347.,-8241.5,-2006.5,-3457.9,-4580.2,-18619.,-298.97,-21550.,-6453.7,-4575.1,-3287.4,94.076,3351.4,3055.9,1579.3,458.97,3114.9,1686.6,0.0000,6685.9,4449.7,4252.8,3658.0,0.0000,-634.64,-215.34,-102.39,-65.309,-115.04,-587.69,0.0000,-1096.2,-1746.6,-756.08,-1462.2
245.0000000000,6255.7,2921.8,3962.8,3063.0,505.16,4098.6,4997.8,858.76,6948.0,2670.8,3466.8,2366.2,0.0000,-10339.,-8239.3,-2006.1,-3454.9,-4573.8,-18612.,-298.30,-21543.,-6454.3,-4575.5,-3286.9,93.792,3341.3,3046.7,1576.7,457.52,3111.5,1686.6,0.0000,6683.8,4449.7,4252.8,3658.0,0.0000,-632.40,-214.53,-102.16,-65.101,-115.01,-587.69,0.0000,-1096.1,-1745.9,-756.15,-1461.4
246.0000000000,6048.2,2922.2,3847.6,2998.1,439.79,4103.3,4962.1,858.77,6956.2,2668.1,3466.7,2351.4,0.0000,-10331.,-8237.0,-2005.7,-3451.9,-4567.4,-18606.,-297.71,-21536.,-6454.9,-4575.8,-3286.5,153.76,3475.6,3111.1,1621.9,466.89,3141.2,1686.6,89.008,6735.5,4471.9,4268.3,3670.9,0.0000,-634.21,-216.20,-102.48,-65.337,-115.64,-587.69,-4.0805,-1096.4,-1745.2,-756.29,-1461.9
247.0000000000,5611.5,2925.3,2843.9,2999.9,411.13,4110.7,4962.4,845.31,6964.6,2667.2,3466.6,2349.6,0.0000,-10323.,-8234.7,-2005.2,-3448.8,-4560.9,-18599.,-297.05,-21530.,-6455.5,-4576.1,-3286.0,93.863,3343.8,3049.0,1580.1,457.90,3119.6,1686.6,0.0000,6688.7,4449.7,4252.8,3658.0,0.0000,-632.24,-214.42,-102.31,-65.130,-115.50,-587.69,0.0000,-1096.1,-1744.5,-756.29,-1460.0
248.0000000000,5579.9,2927.3,2844.5,2996.1,411.38,3978.0,4962.7,836.47,6968.6,2667.9,3458.9,2350.3,0.0000,-10315.,-8232.4,-2004.5,-3445.8,-4554.5,-18592.,-296.44,-21523.,-6456.1,-4576.4,-3285.6,154.14,3351.9,3157.9,1585.6,494.83,3131.3,1686.6,0.0000,6695.8,4449.7,4252.8,3658.0,0.0000,-633.44,-216.97,-102.62,-65.523,-116.04,-587.69,0.0000,-1096.1,-1743.8,-756.36,-1459.3
249.0000000000,5579.9,2932.2,2848.6,2935.4,411.77,3864.9,4928.0,822.90,6971.8,2668.6,3443.2,2351.0,0.0000,-10307.,-8230.2,-2003.9,-3442.8,-4548.1,-18585.,-295.82,-21517.,-6456.7,-4576.7,-3285.1,126.64,3358.0,3104.4,1588.2,484.38,3136.0,1686.6,0.0000,6698.6,4449.7,4252.8,3658.0,0.0000,-634.20,-215.95,-102.79,-65.547,-116.31,-587.69,0.0000,-1096.1,-1743.1,-756.43,-1458.6
250.0000000000,5580.0,2934.8,2850.9,2937.7,412.02,3782.0,4899.6,822.90,6973.7,2659.5,3429.4,2351.7,0.0000,-10299.,-8228.1,-2003.2,-3439.9,-4541.8,-18579.,-295.16,-21510.,-6457.3,-4577.0,-3284.6,94.065,3351.0,3055.6,1586.0,458.92,3132.5,1686.6,0.0000,6696.5,4449.7,4252.8,3658.0,0.0000,-632.63,-214.48,-102.62,-65.238,-116.26,-587.69,0.0000,-1096.1,-1742.4,-756.50,-1458.0
251.0000000000,4864.4,2932.4,2849.8,2938.9,411.67,3760.1,4847.2,815.43,6974.9,2650.2,3413.2,2352.4,0.0000,-10290.,-8225.7,-2002.6,-3436.9,-4535.5,-18572.,-294.50,-21504.,-6457.8,-4577.3,-3284.0,93.814,3342.1,3047.4,1583.4,457.73,3128.6,1686.6,0.0000,6694.2,4449.7,4252.8,3658.0,0.0000,-630.61,-213.78,-102.40,-65.053,-116.20,-587.69,0.0000,-1096.0,-1741.7,-756.57,-1457.3
252.0000000000,4539.7,2929.8,2847.2,2939.4,411.04,3712.5,4836.6,754.20,6910.2,2650.9,3410.7,2353.1,0.0000,-10282.,-8223.2,-2001.8,-3433.8,-4529.2,-18566.,-293.89,-21497.,-6458.4,-4577.6,-3283.5,93.755,3377.8,3045.5,1618.8,457.50,3153.3,1686.6,0.0000,6729.7,4449.7,4263.0,3660.2,0.0000,-629.97,-213.50,-102.45,-65.000,-116.67,-587.69,0.0000,-1096.3,-1741.0,-756.67,-1456.8
253.0000000000,4438.0,2927.1,2843.6,2900.0,410.31,3699.2,4836.9,751.20,6866.8,2651.6,3410.6,2345.2,0.0000,-10273.,-8220.5,-2001.1,-3430.8,-4522.8,-18559.,-293.26,-21491.,-6458.9,-4577.9,-3283.0,93.498,3330.8,3037.1,1583.6,456.28,3132.7,1686.6,0.0000,6696.8,4449.7,4252.8,3658.0,0.0000,-627.82,-212.77,-102.25,-64.810,-116.53,-587.69,0.0000,-1096.0,-1740.4,-756.68,-1455.9
254.0000000000,4437.8,2923.1,2839.2,2871.5,409.70,3649.8,4801.9,751.22,6711.8,2652.3,3410.6,2336.4,0.0000,-10263.,-8217.6,-2000.3,-3427.8,-4516.5,-18552.,-292.65,-21484.,-6459.5,-4578.2,-3282.4,93.399,3327.3,3033.9,1583.7,455.83,3134.0,1686.6,0.0000,6697.6,4449.7,4252.8,3658.0,0.0000,-626.82,-212.40,-102.20,-64.729,-116.66,-587.69,0.0000,-1096.0,-1739.7,-756.73,-1455.3
255.0000000000,4380.2,2919.3,2835.3,2871.8,408.86,3551.6,4766.2,751.23,6689.6,2653.0,3410.5,2322.1,0.0000,-10254.,-8214.6,-1999.5,-3424.7,-4510.2,-18546.,-292.03,-21478.,-6460.0,-4578.5,-3281.8,93.109,3317.0,3024.5,1580.8,454.45,3129.9,1686.6,0.0000,6695.1,4449.7,4252.8,3658.0,0.0000,-624.53,-211.59,-101.95,-64.516,-116.58,-587.69,0.0000,-1095.9,-1739.0,-756.79,-1454.6
256.0000000000,4246.8,2913.5,2828.8,2852.8,407.89,3545.5,4685.4,752.06,6690.3,2643.4,3410.5,2310.6,0.0000,-10244.,-8211.3,-1998.6,-3421.6,-4503.9,-18539.,-291.41,-21471.,-6460.5,-4578.9,-3281.3,92.813,3306.4,3014.9,1577.9,453.04,3125.7,1686.6,0.0000,6692.6,4449.7,4252.8,3658.0,0.0000,-622.21,-210.76,-101.70,-64.297,-116.50,-587.69,0.0000,-1095.8,-1738.3,-756.84,-1454.0
257.0000000000,4112.1,2904.6,2822.2,2803.2,406.72,3545.1,4590.9,714.23,6690.6,2627.2,3410.4,2302.2,0.0000,-10234.,-8207.9,-1997.6,-3418.5,-4497.6,-18533.,-290.80,-21465.,-6461.0,-4579.2,-3280.7,92.517,3295.9,3005.3,1575.0,451.63,3121.3,1686.6,0.0000,6690.1,4449.7,4252.8,3658.0,0.0000,-619.88,-209.93,-101.45,-64.079,-116.40,-587.69,0.0000,-1095.8,-1737.7,-756.89,-1453.3
258.0000000000,3871.1,2883.5,2817.3,2796.3,405.49,3542.9,4463.4,686.16,6690.7,2615.7,3410.3,2302.9,0.0000,-10223.,-8204.2,-1996.6,-3415.4,-4491.2,-18526.,-290.20,-21458.,-6461.5,-4579.6,-3280.1,92.219,3285.2,2995.6,1571.9,450.21,3116.8,1686.6,0.0000,6687.4,4449.7,4252.8,3658.0,0.0000,-617.53,-209.09,-101.19,-63.859,-116.30,-587.69,0.0000,-1095.7,-1737.0,-756.94,-1452.6
259.0000000000,3602.6,2876.2,2810.7,2687.2,404.26,3541.1,4289.2,656.15,6690.9,2616.4,3410.3,2303.6,0.0000,-10212.,-8200.3,-1995.6,-3412.3,-4484.8,-18520.,-289.60,-21452.,-6462.0,-4579.9,-3279.5,91.916,3274.4,2985.8,1568.8,448.76,3112.0,1686.6,0.0000,6684.5,4449.7,4252.8,3658.0,0.0000,-615.14,-208.23,-100.92,-63.635,-116.18,-587.69,0.0000,-1095.7,-1736.3,-756.99,-1452.0
260.0000000000,3227.1,2870.2,2804.2,2621.6,403.35,3539.8,4267.7,630.77,6691.2,2612.4,3410.2,2304.2,0.0000,-10201.,-8196.3,-1994.5,-3409.1,-4478.4,-18513.,-289.03,-21445.,-6462.5,-4580.3,-3278.9,91.878,3273.1,2984.5,1570.1,448.61,3115.8,1686.6,0.0000,6686.8,4449.7,4252.8,3658.0,0.0000,-614.52,-207.97,-100.95,-63.595,-116.39,-587.69,0.0000,-1095.6,-1735.7,-757.04,-1451.3
261.0000000000,3155.0,2868.9,2803.4,2545.7,403.12,3539.1,4248.2,627.16,6691.0,2612.8,3387.7,2304.9,0.0000,-10191.,-8192.4,-1993.4,-3406.0,-4472.0,-18507.,-288.49,-21439.,-6463.1,-4580.6,-3278.4,103.13,3302.4,3011.4,1582.6,456.70,3132.4,1686.6,22.467,6707.4,4458.3,4264.2,3666.1,0.0000,-615.61,-208.70,-101.20,-63.775,-116.83,-587.69,-1.0298,-1095.8,-1735.0,-757.14,-1451.4
262.0000000000,3067.6,2869.1,2803.8,2525.3,403.16,3493.1,4141.5,627.17,6635.8,2613.5,3373.1,2305.5,0.0000,-10180.,-8188.8,-1992.4,-3403.0,-4465.7,-18501.,-287.92,-21432.,-6463.6,-4580.9,-3277.8,91.927,3274.9,2986.1,1572.9,448.89,3122.7,1686.6,0.0000,6691.0,4449.7,4252.8,3658.0,0.0000,-614.14,-207.74,-101.07,-63.604,-116.78,-587.69,0.0000,-1095.6,-1734.3,-757.14,-1450.0
263.0000000000,2950.0,2899.9,2832.3,2493.7,409.46,3474.4,4082.2,627.18,6609.7,2614.2,3373.1,2292.1,0.0000,-10173.,-8186.6,-1991.7,-3400.3,-4459.6,-18494.,-287.60,-21426.,-6464.4,-4581.2,-3277.8,335.35,3899.1,3533.3,1670.9,500.76,3264.3,1686.9,318.47,6800.4,4475.0,4284.1,3682.4,0.0000,-648.09,-227.10,-105.88,-67.239,-121.41,-587.69,-14.597,-1096.7,-1733.7,-757.33,-1451.5
264.0000000000,2896.6,3000.3,2925.3,2499.7,424.59,3519.7,3963.5,616.78,6578.5,2614.8,3373.0,2306.6,0.0000,-10174.,-8189.0,-1995.1,-3398.4,-4456.6,-18488.,-287.26,-21423.,-6465.2,-4581.6,-3277.8,1760.1,5110.9,4930.4,2383.9,623.35,4952.4,1696.5,1224.5,7854.9,4534.9,4370.7,3762.0,0.0000,-689.31,-266.11,-131.06,-71.893,-184.68,-587.86,-56.122,-1108.0,-1733.1,-757.76,-1457.7
265.0000000000,2821.6,3104.8,3026.9,2667.7,446.77,3790.5,3888.3,585.25,6614.4,2606.4,3373.0,2277.5,0.0000,-10182.,-8195.1,-2003.3,-3397.1,-4461.4,-18482.,-286.66,-21425.,-6465.7,-4581.9,-3277.0,104.66,3728.5,3399.8,2387.8,715.17,4890.2,1692.4,0.0000,7917.6,4479.0,4295.6,3792.9,0.0000,-698.77,-236.49,-132.32,-73.787,-184.67,-587.79,0.0000,-1108.5,-1732.5,-757.48,-1459.7
266.0000000000,2692.2,3107.2,3088.2,2826.4,462.45,4048.1,3845.3,550.54,6677.8,2596.3,3373.1,2266.4,0.0000,-10192.,-8201.4,-2014.2,-3395.9,-4476.0,-18476.,-285.98,-21430.,-6466.0,-4582.2,-3276.0,104.79,3733.0,3403.8,2307.9,539.45,4870.4,1691.9,0.0000,7753.2,4462.8,4272.4,3676.1,0.0000,-699.62,-236.87,-132.40,-72.678,-184.99,-587.78,0.0000,-1107.0,-1731.9,-757.42,-1449.3
267.0000000000,2671.3,3109.6,3112.4,2934.2,465.31,4200.5,3825.0,519.44,6741.8,2581.2,3373.0,2267.1,0.0000,-10200.,-8206.5,-2024.6,-3394.3,-4487.9,-18469.,-285.33,-21445.,-6466.3,-4582.5,-3275.1,104.64,3727.6,3398.9,2298.5,526.74,4859.2,1691.4,0.0000,7744.9,4453.8,4259.5,3664.4,0.0000,-698.65,-236.62,-132.30,-72.500,-185.41,-587.77,0.0000,-1106.9,-1731.2,-757.41,-1447.6
268.0000000000,2648.3,3117.1,3121.5,2892.7,465.04,4297.4,3825.2,518.69,6750.1,2578.0,3372.8,2260.0,0.0000,-10206.,-8210.5,-2035.7,-3392.6,-4495.8,-18463.,-284.71,-21465.,-6466.6,-4582.7,-3274.2,104.36,3717.7,3389.9,2293.8,519.87,4854.6,1691.0,0.0000,7741.5,4450.5,4254.2,3659.3,0.0000,-696.83,-236.08,-132.12,-72.274,-185.89,-587.77,0.0000,-1106.8,-1730.6,-757.44,-1446.6
269.0000000000,2534.8,3096.6,3129.4,2892.1,464.00,4373.0,3825.5,488.60,6868.0,2578.6,3372.8,2250.9,0.0000,-10211.,-8213.5,-2047.4,-3390.6,-4501.3,-18457.,-284.11,-21478.,-6467.0,-4583.0,-3273.4,104.03,3705.8,3379.1,2291.6,516.85,4853.4,1690.3,0.0000,7740.9,4449.7,4252.9,3658.1,0.0000,-694.62,-235.40,-131.90,-72.034,-186.38,-587.75,0.0000,-1106.8,-1729.9,-757.48,-1445.9
270.0000000000,2297.9,3051.8,3131.0,2873.4,462.69,4541.0,3825.6,454.72,6999.8,2578.0,3372.9,2234.2,0.0000,-10215.,-8215.6,-2055.7,-3388.5,-4505.3,-18451.,-283.54,-21486.,-6467.4,-4583.3,-3272.7,103.66,3692.8,3367.3,2289.9,515.02,4853.1,1690.3,0.0000,7740.9,4449.7,4252.8,3658.0,0.0000,-692.18,-234.63,-131.65,-71.779,-186.86,-587.75,0.0000,-1106.8,-1729.3,-757.52,-1445.2
271.0000000000,2173.3,3049.5,3124.1,2882.5,461.23,4702.7,3803.9,437.49,7110.7,2574.8,3372.8,2215.7,0.0000,-10217.,-8217.0,-2062.1,-3386.4,-4508.3,-18445.,-282.97,-21493.,-6467.8,-4583.6,-3271.9,103.28,3679.2,3354.8,2288.2,513.23,4853.0,1689.8,0.0000,7740.9,4449.7,4252.8,3658.0,0.0000,-689.58,-233.80,-131.40,-71.509,-187.34,-587.75,0.0000,-1106.7,-1728.6,-757.57,-1444.6
272.0000000000,2111.7,3049.7,3122.7,2898.3,460.42,4755.4,3602.0,411.24,7154.7,2575.5,3372.7,2196.0,0.0000,-10218.,-8218.3,-2067.5,-3384.1,-4510.8,-18440.,-282.44,-21499.,-6468.2,-4583.8,-3271.3,168.17,3825.2,3425.5,2290.9,584.84,4872.4,1689.8,0.0000,7740.9,4449.7,4339.2,3748.9,0.0000,-690.94,-235.60,-131.51,-72.103,-187.94,-587.74,0.0000,-1106.7,-1728.0,-758.00,-1451.6
273.0000000000,2035.6,3050.4,3123.9,2904.0,459.80,4774.4,3508.4,374.95,7177.9,2576.1,3372.6,2158.5,0.0000,-10218.,-8219.3,-2072.2,-3381.9,-4513.0,-18434.,-281.88,-21505.,-6468.6,-4584.1,-3270.5,103.14,3674.5,3350.5,2287.6,512.61,4853.0,1689.4,0.0000,7740.9,4449.7,4252.8,3658.0,0.0000,-688.58,-233.55,-131.31,-71.407,-188.27,-587.74,0.0000,-1106.7,-1727.4,-757.66,-1443.3
274.0000000000,2060.6,3046.2,3120.9,2910.5,458.99,4776.9,3508.6,348.55,7182.4,2576.8,3372.5,2128.9,0.0000,-10217.,-8220.0,-2076.5,-3379.6,-4514.9,-18428.,-281.33,-21510.,-6469.0,-4584.4,-3269.8,102.78,3661.4,3338.6,2286.0,510.90,4852.8,1689.2,0.0000,7740.9,4449.7,4252.8,3658.0,0.0000,-686.04,-232.72,-131.07,-71.146,-188.72,-587.73,0.0000,-1106.6,-1726.7,-757.70,-1442.7
275.0000000000,2003.4,3039.0,3116.1,2893.7,457.69,4787.8,3508.7,332.00,7162.7,2573.5,3372.6,2128.6,0.0000,-10215.,-8220.2,-2080.4,-3377.3,-4516.7,-18422.,-280.77,-21515.,-6469.4,-4584.6,-3269.0,102.39,3647.5,3325.9,2284.2,509.08,4852.7,1689.2,0.0000,7740.9,4449.7,4252.8,3658.0,0.0000,-683.32,-231.83,-130.81,-70.868,-189.16,-587.73,0.0000,-1106.6,-1726.1,-757.75,-1442.1
276.0000000000,1910.6,3032.6,3106.4,2839.9,456.21,4812.2,3508.9,319.90,7145.8,2570.5,3372.7,2129.2,0.0000,-10213.,-8219.9,-2084.0,-3374.9,-4518.9,-18417.,-280.22,-21520.,-6469.8,-4584.9,-3268.3,101.99,3633.3,3313.0,2282.4,507.23,4852.6,1689.0,0.0000,7740.9,4449.7,4252.8,3658.0,0.0000,-680.53,-230.90,-130.54,-70.583,-189.58,-587.73,0.0000,-1106.6,-1725.4,-757.79,-1441.5
277.0000000000,1868.1,3022.7,3096.0,2851.2,454.59,4762.8,3497.2,287.18,7149.8,2552.2,3361.3,2130.1,0.0000,-10209.,-8219.1,-2087.3,-3372.5,-4521.0,-18411.,-279.68,-21525.,-6470.2,-4585.2,-3267.5,101.59,3619.0,3299.9,2280.6,505.34,4852.4,1688.8,0.0000,7740.9,4449.7,4252.8,3658.0,0.0000,-677.68,-229.95,-130.27,-70.294,-189.98,-587.73,0.0000,-1106.5,-1724.8,-757.84,-1440.9
278.0000000000,1795.8,3012.0,3084.9,2850.5,452.81,4776.0,3445.9,277.95,7146.5,2545.9,3353.9,2127.6,0.0000,-10205.,-8217.9,-2090.3,-3370.0,-4523.2,-18406.,-279.14,-21529.,-6470.6,-4585.4,-3266.8,101.19,3604.7,3286.9,2278.8,503.47,4852.3,1687.6,0.0000,7740.9,4449.7,4252.8,3658.0,0.0000,-674.83,-228.98,-130.00,-70.006,-190.39,-587.70,0.0000,-1106.5,-1724.2,-757.88,-1440.3
279.0000000000,1717.1,3003.0,3074.0,2849.7,451.32,4777.7,3446.0,268.72,7086.5,2536.7,3353.9,2108.6,0.0000,-10200.,-8216.2,-2093.1,-3367.5,-4525.2,-18400.,-278.60,-21534.,-6471.0,-4585.7,-3266.0,100.87,3593.5,3276.7,2277.4,502.01,4852.2,1686.8,0.0000,7740.9,4449.7,4252.8,3658.0,0.0000,-672.55,-228.21,-129.79,-69.778,-190.81,-587.69,0.0000,-1106.5,-1723.5,-757.92,-1439.7
280.0000000000,1698.2,2994.9,3065.4,2849.7,449.96,4779.3,3446.2,259.53,7037.0,2526.7,3354.0,2095.8,0.0000,-10194.,-8214.3,-2095.7,-3364.9,-4527.0,-18395.,-278.07,-21538.,-6471.4,-4585.9,-3265.3,100.56,3582.3,3266.4,2276.0,500.54,4852.1,1686.7,0.0000,7740.9,4449.7,4252.8,3658.0,0.0000,-670.23,-227.41,-129.58,-69.548,-191.21,-587.69,0.0000,-1106.5,-1722.9,-757.97,-1439.1
281.0000000000,1599.6,2986.2,3060.0,2848.6,448.61,4791.8,3386.6,242.66,7049.4,2527.3,3354.0,2096.3,0.0000,-10188.,-8212.1,-2098.1,-3362.3,-4529.0,-18389.,-277.55,-21541.,-6471.8,-4586.2,-3264.5,100.23,3570.6,3255.8,2274.6,499.01,4852.0,1686.6,0.0000,7740.9,4449.7,4252.8,3658.0,0.0000,-667.82,-226.58,-129.37,-69.310,-191.61,-587.69,0.0000,-1106.4,-1722.3,-758.01,-1438.6
282.0000000000,1589.8,2978.8,3056.0,2815.3,447.28,4770.2,3327.0,217.74,7054.3,2528.0,3354.0,2092.7,0.0000,-10182.,-8209.5,-2100.4,-3359.7,-4531.0,-18384.,-277.04,-21545.,-6472.2,-4586.4,-3263.8,99.895,3558.7,3244.9,2273.1,497.45,4851.9,1686.6,0.0000,7740.9,4449.7,4252.8,3658.0,0.0000,-665.36,-225.73,-129.14,-69.068,-192.00,-587.69,0.0000,-1106.4,-1721.7,-758.05,-1438.0
283.0000000000,1589.4,2969.8,3047.0,2779.0,445.95,4742.7,3192.8,205.89,7062.1,2528.6,3354.0,2079.2,0.0000,-10175.,-8206.8,-2102.5,-3357.1,-4532.8,-18379.,-276.53,-21548.,-6472.6,-4586.7,-3263.0,99.557,3546.7,3234.0,2271.6,495.87,4851.8,1686.6,0.0000,7740.9,4449.7,4252.8,3658.0,0.0000,-662.86,-224.85,-128.92,-68.822,-192.38,-587.69,0.0000,-1106.4,-1721.0,-758.10,-1437.5
284.0000000000,1437.3,2960.5,3041.2,2778.9,444.56,4745.1,3129.4,203.32,7085.5,2529.3,3354.1,2079.8,0.0000,-10168.,-8203.8,-2104.5,-3354.4,-4534.3,-18374.,-276.02,-21551.,-6473.0,-4586.9,-3262.3,99.195,3533.8,3222.2,2269.9,494.18,4851.6,1686.6,0.0000,7740.9,4449.7,4252.8,3658.0,0.0000,-660.18,-223.92,-128.68,-68.559,-192.75,-587.69,0.0000,-1106.3,-1720.4,-758.14,-1436.9
285.0000000000,1257.5,2950.6,3033.4,2777.7,443.13,4739.5,2997.8,206.19,7094.4,2530.0,3354.1,2080.4,0.0000,-10161.,-8200.6,-2106.3,-3351.7,-4535.5,-18368.,-275.51,-21554.,-6473.4,-4587.2,-3261.5,98.832,3520.8,3210.4,2268.3,492.49,4851.5,1686.6,0.0000,7740.9,4449.7,4252.8,3658.0,0.0000,-657.49,-222.97,-128.43,-68.296,-193.12,-587.69,0.0000,-1106.3,-1719.7,-758.18,-1436.4
286.0000000000,1131.8,2940.2,3023.2,2776.5,441.71,4674.3,2913.3,205.32,7101.8,2530.6,3353.9,2073.8,0.0000,-10153.,-8197.2,-2108.1,-3349.0,-4536.5,-18363.,-275.00,-21557.,-6473.8,-4587.4,-3260.7,98.488,3508.6,3199.2,2266.8,490.88,4851.4,1686.6,0.0000,7740.9,4449.7,4252.8,3658.0,0.0000,-654.92,-222.06,-128.21,-68.046,-193.49,-587.69,0.0000,-1106.3,-1719.1,-758.22,-1435.8
287.0000000000,1010.2,2933.0,3015.1,2775.2,440.76,4673.9,2875.2,184.05,7105.8,2531.3,3353.7,2063.3,0.0000,-10145.,-8193.6,-2109.7,-3346.3,-4537.7,-18358.,-274.51,-21559.,-6474.2,-4587.7,-3260.0,106.90,3509.1,3199.7,2266.8,492.20,4855.3,1686.6,5.4900,7742.4,4450.6,4262.0,3665.5,0.0000,-654.72,-221.96,-128.21,-68.052,-193.87,-587.69,-0.25156,-1106.3,-1718.5,-758.31,-1435.9
288.0000000000,957.03,2932.8,3013.8,2770.6,440.90,4656.7,2864.6,166.72,7105.8,2531.9,3353.5,2063.9,0.0000,-10137.,-8190.3,-2111.2,-3343.6,-4539.4,-18353.,-274.04,-21562.,-6474.7,-4587.9,-3259.3,187.83,3606.8,3373.0,2283.5,530.38,4877.8,1686.6,98.355,7767.8,4466.6,4291.5,3697.8,0.0000,-657.29,-226.16,-128.48,-68.567,-194.37,-587.69,-4.5066,-1106.5,-1717.9,-758.48,-1438.0
289.0000000000,957.56,2956.8,3036.0,2706.1,445.45,4573.3,2812.0,160.24,7105.6,2532.5,3353.3,2064.5,0.0000,-10132.,-8188.3,-2112.9,-3341.2,-4540.6,-18348.,-273.66,-21564.,-6475.2,-4588.1,-3258.9,742.98,4136.5,4172.2,2324.2,588.95,4915.2,1686.6,599.11,7807.5,4498.5,4334.7,3741.4,0.0000,-678.02,-247.83,-130.49,-70.951,-194.96,-587.69,-27.451,-1106.9,-1717.3,-758.71,-1441.1
290.0000000000,924.74,2999.8,3076.9,2659.1,451.50,4553.7,2812.1,148.90,7105.6,2533.1,3353.2,2065.0,0.0000,-10130.,-8188.4,-2114.6,-3339.2,-4541.3,-18343.,-273.17,-21566.,-6475.6,-4588.4,-3258.1,102.77,3661.2,3338.4,2286.1,527.76,4853.8,1686.6,0.0000,7741.5,4451.9,4256.8,3663.6,0.0000,-682.39,-231.31,-131.06,-71.095,-194.89,-587.69,0.0000,-1106.2,-1716.6,-758.41,-1434.2
291.0000000000,798.46,3021.2,3099.4,2577.9,456.05,4571.1,2812.2,124.79,7105.6,2533.7,3353.3,2061.0,0.0000,-10129.,-8188.7,-2116.2,-3337.1,-4541.8,-18338.,-272.64,-21568.,-6476.0,-4588.6,-3257.2,102.81,3662.4,3339.5,2286.2,523.36,4853.5,1686.6,0.0000,7741.3,4451.3,4255.0,3661.0,0.0000,-682.46,-231.35,-131.08,-71.087,-195.22,-587.69,0.0000,-1106.2,-1716.0,-758.44,-1433.5
292.0000000000,663.69,3027.8,3108.4,2579.4,457.18,4571.0,2812.3,93.584,7094.6,2534.3,3353.4,2048.1,0.0000,-10128.,-8188.7,-2117.8,-3335.0,-4542.0,-18333.,-272.10,-21570.,-6476.3,-4588.9,-3256.3,102.70,3658.6,3336.1,2285.6,515.71,4853.0,1686.6,0.0000,7740.9,4450.2,4253.4,3658.9,0.0000,-681.60,-231.07,-131.01,-70.963,-195.55,-587.69,0.0000,-1106.1,-1715.4,-758.47,-1432.8
293.0000000000,581.36,3029.5,3110.6,2520.9,456.88,4578.2,2797.2,77.036,7095.0,2535.2,3353.3,2048.6,0.0000,-10126.,-8188.3,-2119.2,-3332.8,-4542.0,-18328.,-271.58,-21573.,-6476.6,-4589.1,-3255.5,102.52,3652.2,3330.2,2284.8,511.56,4852.8,1686.6,0.0000,7740.9,4449.8,4252.9,3658.2,0.0000,-680.25,-230.62,-130.89,-70.811,-195.87,-587.69,0.0000,-1106.1,-1714.8,-758.51,-1432.2
294.0000000000,583.50,3027.5,3112.1,2494.8,456.13,4528.8,2685.0,75.024,7099.8,2535.9,3353.1,2049.2,0.0000,-10123.,-8187.6,-2120.5,-3330.5,-4541.8,-18323.,-271.06,-21575.,-6477.0,-4589.3,-3254.6,102.29,3643.9,3322.6,2283.8,509.21,4852.7,1686.6,0.0000,7740.9,4449.7,4252.8,3658.0,0.0000,-678.53,-230.04,-130.74,-70.636,-196.19,-587.69,0.0000,-1106.1,-1714.1,-758.55,-1431.6
295.0000000000,583.31,3024.9,3109.4,2494.6,455.18,4518.7,2629.5,79.071,7102.9,2536.5,3353.0,2049.6,0.0000,-10120.,-8186.5,-2121.7,-3328.2,-4541.5,-18318.,-270.56,-21578.,-6477.3,-4589.6,-3253.8,102.03,3634.8,3314.4,2282.6,507.55,4852.6,1686.6,0.0000,7740.9,4449.7,4252.8,3658.0,0.0000,-676.67,-229.41,-130.57,-70.450,-196.51,-587.69,0.0000,-1106.1,-1713.5,-758.59,-1431.1
296.0000000000,583.04,2994.5,3103.0,2495.3,454.16,4511.9,2585.2,61.860,7105.1,2537.1,3352.9,2050.1,0.0000,-10117.,-8185.0,-2122.9,-3325.8,-4541.0,-18313.,-270.05,-21580.,-6477.7,-4589.8,-3253.0,101.77,3625.5,3305.9,2281.5,506.22,4852.5,1686.6,0.0000,7740.9,4449.7,4252.8,3658.0,0.0000,-674.76,-228.76,-130.39,-70.261,-196.82,-587.69,0.0000,-1106.0,-1712.9,-758.63,-1430.6
297.0000000000,582.74,2946.4,3096.5,2495.0,453.09,4502.1,2513.8,58.316,7106.4,2537.7,3352.8,2035.8,0.0000,-10112.,-8183.3,-2124.0,-3323.4,-4540.4,-18308.,-269.56,-21582.,-6478.0,-4590.0,-3252.2,101.49,3615.6,3296.8,2280.2,504.90,4852.4,1686.6,0.0000,7740.9,4449.7,4252.8,3658.0,0.0000,-672.70,-228.06,-130.21,-70.059,-197.12,-587.69,0.0000,-1106.0,-1712.3,-758.67,-1430.0
298.0000000000,537.06,2941.5,3090.3,2494.1,451.98,4489.4,2494.7,52.156,7116.6,2538.4,3352.8,2033.3,0.0000,-10107.,-8181.3,-2125.0,-3320.9,-4539.7,-18303.,-269.06,-21584.,-6478.3,-4590.2,-3251.4,101.20,3605.2,3287.3,2278.9,503.54,4852.3,1686.6,0.0000,7740.9,4449.7,4252.8,3658.0,0.0000,-670.56,-227.32,-130.01,-69.849,-197.43,-587.69,0.0000,-1106.0,-1711.6,-758.71,-1429.5
299.0000000000,474.12,2935.9,3083.1,2493.0,450.82,4483.2,2494.8,40.782,7121.5,2539.0,3352.8,2033.9,0.0000,-10101.,-8179.1,-2126.0,-3318.4,-4538.8,-18298.,-268.56,-21585.,-6478.7,-4590.5,-3250.6,100.90,3594.5,3277.6,2277.6,502.14,4852.2,1686.6,0.0000,7740.9,4449.7,4252.8,3658.0,0.0000,-668.35,-226.56,-129.81,-69.632,-197.72,-587.69,0.0000,-1106.0,-1711.0,-758.75,-1429.0
300.0000000000,376.51,2928.5,3076.6,2491.9,449.62,4482.8,2481.8,40.785,7067.9,2539.6,3352.8,2034.3,0.0000,-10095.,-8176.7,-2126.9,-3315.9,-4537.9,-18293.,-268.07,-21587.,-6479.0,-4590.7,-3249.8,100.59,3583.4,3267.5,2276.2,500.69,4852.1,1686.6,0.0000,7740.9,4449.7,4252.8,3658.0,0.0000,-666.06,-225.76,-129.61,-69.407,-198.02,-587.69,0.0000,-1105.9,-1710.4,-758.78,-1428.5
301.0000000000,325.76,2921.3,3068.1,2490.8,448.39,4470.0,2368.3,25.024,7038.1,2540.2,3352.7,2034.7,0.0000,-10088.,-8174.2,-2127.7,-3313.3,-4536.9,-18288.,-267.58,-21588.,-6479.3,-4590.9,-3249.0,100.28,3572.3,3257.4,2274.8,499.23,4852.0,1686.6,0.0000,7740.9,4449.7,4252.8,3658.0,0.0000,-663.75,-224.96,-129.40,-69.181,-198.30,-587.69,0.0000,-1105.9,-1709.8,-758.82,-1427.9
302.0000000000,325.43,2913.1,3059.0,2493.8,447.13,4464.1,2309.8,22.967,6986.4,2540.8,3352.6,2022.6,0.0000,-10081.,-8171.4,-2128.5,-3310.7,-4535.8,-18283.,-267.09,-21589.,-6479.7,-4591.1,-3248.1,99.951,3560.7,3246.8,2273.3,497.71,4851.9,1686.6,0.0000,7740.9,4449.7,4252.8,3658.0,0.0000,-661.34,-224.11,-129.18,-68.945,-198.59,-587.69,0.0000,-1105.9,-1709.1,-758.86,-1427.4
303.0000000000,325.09,2904.1,3048.8,2461.2,445.84,4463.6,2261.1,22.970,6986.5,2541.4,3352.6,2008.3,0.0000,-10074.,-8168.4,-2129.2,-3308.1,-4534.6,-18278.,-266.60,-21590.,-6480.0,-4591.4,-3247.3,99.624,3549.0,3236.1,2271.9,496.18,4851.8,1686.6,0.0000,7740.9,4449.7,4252.8,3658.0,0.0000,-658.91,-223.26,-128.96,-68.708,-198.87,-587.69,0.0000,-1105.9,-1708.6,-758.90,-1426.9
304.0000000000,324.75,2895.8,3039.2,2410.5,444.56,4463.2,2238.2,22.973,6956.0,2541.9,3352.6,2000.5,0.0000,-10066.,-8165.3,-2129.9,-3305.5,-4533.3,-18273.,-266.11,-21591.,-6480.3,-4591.6,-3246.4,99.325,3538.4,3226.4,2270.5,494.79,4851.7,1686.6,0.0000,7740.9,4449.7,4252.8,3658.0,0.0000,-656.66,-222.47,-128.76,-68.491,-199.15,-587.69,0.0000,-1105.8,-1708.0,-758.93,-1426.4
305.0000000000,324.44,2887.9,3030.8,2357.5,443.36,4462.6,2119.0,23.637,6915.1,2542.5,3352.5,2001.1,0.0000,-10057.,-8162.0,-2130.5,-3302.9,-4532.0,-18268.,-265.63,-21592.,-6480.6,-4591.8,-3245.6,99.045,3528.4,3217.3,2269.3,493.48,4851.6,1686.6,0.0000,7740.9,4449.7,4252.8,3658.0,0.0000,-654.53,-221.71,-128.58,-68.286,-199.42,-587.69,0.0000,-1105.8,-1707.4,-758.97,-1425.9
306.0000000000,324.16,2880.0,3023.6,2361.5,442.23,4462.1,2114.7,24.564,6914.6,2543.1,3352.6,2001.6,0.0000,-10049.,-8158.6,-2131.2,-3300.2,-4530.6,-18264.,-265.14,-21592.,-6480.9,-4592.1,-3244.8,98.768,3518.6,3208.4,2268.0,492.19,4851.5,1686.6,0.0000,7740.9,4449.7,4252.8,3658.0,0.0000,-652.41,-220.95,-128.39,-68.083,-199.68,-587.69,0.0000,-1105.8,-1706.8,-759.01,-1425.4
307.0000000000,300.44,2872.3,3016.3,2360.9,441.13,4461.8,2084.7,23.479,6914.5,2543.6,3352.6,2002.1,0.0000,-10040.,-8154.9,-2131.7,-3297.6,-4529.1,-18259.,-264.66,-21593.,-6481.2,-4592.3,-3243.9,98.503,3509.1,3199.7,2266.8,490.95,4851.4,1686.6,0.0000,7740.9,4449.7,4252.8,3658.0,0.0000,-650.36,-220.21,-128.22,-67.888,-199.95,-587.69,0.0000,-1105.8,-1706.2,-759.05,-1424.8
308.0000000000,260.62,2867.0,3010.3,2360.1,440.44,4461.4,2051.9,22.728,6914.6,2544.2,3352.5,1985.8,0.0000,-10032.,-8151.2,-2132.3,-3294.9,-4527.5,-18254.,-264.18,-21593.,-6481.5,-4592.5,-3243.1,98.528,3510.0,3200.6,2267.0,491.07,4851.4,1686.6,0.0000,7740.9,4449.7,4252.8,3658.0,0.0000,-650.23,-220.13,-128.23,-67.894,-200.21,-587.69,0.0000,-1105.7,-1705.6,-759.08,-1424.3
309.0000000000,260.35,2863.5,3007.6,2335.0,439.89,4461.0,2052.0,23.541,6914.6,2544.8,3352.5,1985.0,0.0000,-10023.,-8147.7,-2132.8,-3292.3,-4525.9,-18249.,-263.70,-21594.,-6481.8,-4592.8,-3242.2,98.326,3502.8,3194.0,2266.0,490.13,4851.4,1686.6,0.0000,7740.9,4449.7,4252.8,3658.0,0.0000,-648.59,-219.53,-128.10,-67.744,-200.46,-587.69,0.0000,-1105.7,-1705.1,-759.12,-1423.8
310.0000000000,260.03,2858.9,3004.8,2289.1,439.47,4466.4,2023.6,24.317,6914.5,2545.3,3352.3,1985.5,0.0000,-10015.,-8144.4,-2133.3,-3289.6,-4524.2,-18244.,-263.23,-21594.,-6482.1,-4593.0,-3241.4,98.219,3499.0,3190.5,2265.6,489.63,4851.3,1686.6,0.0000,7740.9,4449.7,4252.8,3658.0,0.0000,-647.59,-219.15,-128.03,-67.659,-200.71,-587.69,0.0000,-1105.7,-1704.5,-759.16,-1423.3
311.0000000000,259.92,2855.0,3001.9,2288.4,438.99,4466.0,1967.6,24.319,6914.4,2545.9,3352.2,1986.0,0.0000,-10006.,-8141.1,-2133.8,-3287.0,-4522.5,-18240.,-262.75,-21594.,-6482.4,-4593.3,-3240.5,98.133,3495.9,3187.7,2265.2,489.23,4851.3,1686.6,4.5019,7740.9,4451.5,4252.8,3658.0,0.0000,-646.71,-218.81,-127.97,-67.589,-200.96,-587.69,-0.20622,-1105.7,-1703.9,-759.19,-1422.8
312.0000000000,259.77,2851.1,2997.0,2287.8,438.41,4465.7,1925.1,13.886,6914.4,2546.5,3352.1,1980.7,0.0000,-9998.0,-8137.7,-2134.2,-3284.4,-4520.7,-18235.,-262.28,-21595.,-6482.6,-4593.5,-3239.6,97.894,3487.4,3180.0,2264.1,488.11,4851.2,1686.6,0.0000,7740.9,4449.7,4252.8,3658.0,0.0000,-644.84,-218.13,-127.81,-67.414,-201.20,-587.69,0.0000,-1105.7,-1703.3,-759.23,-1422.3
313.0000000000,259.59,2847.0,2991.9,2287.0,437.91,4465.4,1925.1,5.0396,6911.2,2547.2,3351.9,1969.2,0.0000,-9989.4,-8134.3,-2134.7,-3281.8,-4518.9,-18230.,-261.80,-21595.,-6482.9,-4593.8,-3238.7,97.867,3486.5,3179.1,2264.0,487.99,4851.2,1686.6,0.0000,7740.9,4449.7,4252.8,3658.0,0.0000,-644.36,-217.93,-127.79,-67.385,-201.44,-587.69,0.0000,-1105.6,-1702.8,-759.26,-1421.8
314.0000000000,259.47,2843.4,2987.8,2286.4,437.28,4465.2,1908.0,4.7241,6912.9,2547.7,3351.9,1969.7,0.0000,-9980.9,-8130.8,-2135.1,-3279.1,-4517.0,-18225.,-261.32,-21595.,-6483.2,-4594.0,-3237.8,97.614,3477.5,3170.9,2262.9,486.81,4851.1,1686.6,0.0000,7740.9,4449.7,4252.8,3658.0,0.0000,-642.39,-217.21,-127.62,-67.200,-201.67,-587.69,0.0000,-1105.6,-1702.2,-759.30,-1421.3
315.0000000000,259.25,2837.7,2981.7,2285.9,436.50,4465.1,1861.9,4.7255,6851.9,2548.3,3351.9,1970.3,0.0000,-9972.1,-8127.2,-2135.4,-3276.5,-4515.1,-18221.,-260.84,-21595.,-6483.4,-4594.2,-3236.9,97.358,3468.3,3162.5,2261.7,485.61,4851.0,1686.6,0.0000,7740.9,4449.7,4252.8,3658.0,0.0000,-640.39,-216.49,-127.45,-67.012,-201.90,-587.69,0.0000,-1105.6,-1701.6,-759.33,-1420.8
316.0000000000,259.02,2831.8,2975.1,2287.0,435.52,4464.7,1861.9,4.7268,6848.1,2548.8,3351.8,1970.8,0.0000,-9963.0,-8123.6,-2135.7,-3273.8,-4513.1,-18216.,-260.37,-21595.,-6483.7,-4594.5,-3236.0,97.127,3460.1,3155.0,2260.7,484.53,4851.0,1686.6,0.0000,7740.9,4449.7,4252.8,3658.0,0.0000,-638.56,-215.83,-127.30,-66.842,-202.13,-587.69,0.0000,-1105.6,-1701.1,-759.35,-1420.3
317.0000000000,201.12,2826.5,2968.7,2252.4,434.61,4464.3,1862.0,4.7281,6848.0,2549.3,3351.8,1971.3,0.0000,-9953.8,-8119.8,-2136.0,-3271.2,-4511.1,-18211.,-259.89,-21595.,-6483.9,-4594.7,-3235.1,96.927,3453.0,3148.5,2259.8,483.60,4850.9,1686.6,0.0000,7740.9,4449.7,4252.8,3658.0,0.0000,-636.94,-215.23,-127.16,-66.693,-202.35,-587.69,0.0000,-1105.5,-1700.5,-759.36,-1419.8
318.0000000000,194.67,2820.8,2962.5,2221.1,433.78,4464.0,1801.0,4.7294,6848.1,2549.8,3351.8,1971.8,0.0000,-9944.5,-8116.1,-2136.3,-3268.5,-4509.0,-18206.,-259.42,-21594.,-6484.2,-4594.9,-3234.2,96.730,3445.9,3142.1,2258.9,482.68,4850.8,1686.6,0.0000,7740.9,4449.7,4252.8,3658.0,0.0000,-635.33,-214.63,-127.03,-66.546,-202.57,-587.69,0.0000,-1105.5,-1699.9,-759.37,-1419.4
319.0000000000,194.45,2815.4,2957.0,2220.3,433.01,4407.3,1671.9,4.7307,6848.1,2550.4,3351.8,1972.2,0.0000,-9935.1,-8112.3,-2136.6,-3265.8,-4506.9,-18202.,-258.95,-21594.,-6484.4,-4595.2,-3233.3,96.520,3438.5,3135.3,2258.0,481.70,4850.7,1686.6,0.0000,7740.9,4449.7,4252.8,3658.0,0.0000,-633.63,-214.01,-126.89,-66.391,-202.79,-587.69,0.0000,-1105.5,-1699.4,-759.39,-1418.9
320.0000000000,194.22,2809.3,2951.1,2219.5,432.21,4392.2,1671.9,5.7513,6848.1,2551.0,3351.8,1972.8,0.0000,-9925.6,-8108.4,-2136.8,-3263.1,-4504.8,-18197.,-258.48,-21594.,-6484.6,-4595.4,-3232.5,96.281,3430.0,3127.5,2256.9,480.58,4850.7,1686.6,0.0000,7740.9,4449.7,4252.8,3658.0,0.0000,-631.74,-213.32,-126.73,-66.214,-203.00,-587.69,0.0000,-1105.5,-1698.8,-759.40,-1418.4
321.0000000000,193.97,2802.9,2943.6,2218.6,431.21,4399.5,1622.8,6.3320,6848.1,2551.6,3351.7,1973.3,0.0000,-9915.9,-8104.3,-2137.0,-3260.4,-4502.8,-18192.,-258.00,-21594.,-6484.8,-4595.6,-3231.6,96.024,3420.8,3119.2,2255.8,479.39,4850.6,1686.6,0.0000,7740.9,4449.7,4252.8,3658.0,0.0000,-629.73,-212.59,-126.56,-66.026,-203.14,-587.69,0.0000,-1105.5,-1698.2,-759.41,-1417.9
322.0000000000,193.74,2796.3,2935.9,2217.7,430.20,4402.8,1608.6,6.3333,6848.1,2552.2,3351.6,1973.8,0.0000,-9906.1,-8100.2,-2137.1,-3257.7,-4502.1,-18188.,-257.54,-21593.,-6485.1,-4595.8,-3230.7,95.766,3411.6,3110.8,2254.6,478.18,4850.5,1686.6,0.0000,7740.9,4449.7,4252.8,3658.0,0.0000,-627.71,-211.86,-126.39,-65.837,-203.28,-587.69,0.0000,-1105.4,-1697.7,-759.42,-1417.4
323.0000000000,193.63,2790.4,2929.1,2216.7,429.20,4406.2,1608.7,4.8770,6848.0,2552.7,3351.6,1974.3,0.0000,-9896.1,-8096.1,-2137.3,-3255.0,-4502.8,-18183.,-257.07,-21593.,-6485.3,-4596.0,-3229.8,95.522,3402.9,3102.9,2253.5,477.04,4850.4,1686.6,0.0000,7740.9,4449.7,4252.8,3658.0,0.0000,-625.78,-211.15,-126.23,-65.658,-203.41,-587.69,0.0000,-1105.4,-1697.1,-759.43,-1416.9
324.0000000000,193.37,2783.7,2923.1,2215.7,428.18,4405.8,1608.7,4.5130,6781.9,2553.2,3351.6,1974.8,0.0000,-9885.9,-8092.0,-2137.4,-3252.3,-4504.3,-18178.,-256.60,-21592.,-6485.5,-4596.2,-3229.0,95.268,3393.9,3094.7,2252.4,475.86,4850.3,1686.6,0.0000,7740.9,4449.7,4252.8,3658.0,0.0000,-623.79,-210.42,-126.06,-65.471,-203.53,-587.69,0.0000,-1105.4,-1696.6,-759.44,-1416.4
325.0000000000,193.10,2777.3,2916.7,2214.7,427.14,4405.5,1575.5,4.5142,6780.0,2553.7,3351.6,1975.2,0.0000,-9875.6,-8087.8,-2137.5,-3249.6,-4506.1,-18174.,-256.14,-21592.,-6485.7,-4596.3,-3228.1,95.022,3385.1,3086.7,2251.3,474.71,4850.2,1686.6,0.0000,7740.9,4449.7,4252.8,3658.0,0.0000,-621.84,-209.71,-125.89,-65.290,-203.64,-587.69,0.0000,-1105.4,-1696.0,-759.45,-1415.9
326.0000000000,192.98,2771.3,2912.0,2208.2,426.34,4408.3,1545.4,4.5155,6780.1,2554.3,3351.6,1975.8,0.0000,-9865.3,-8083.7,-2137.6,-3246.9,-4507.9,-18169.,-255.67,-21591.,-6485.9,-4596.5,-3227.2,94.919,3381.5,3083.3,2250.8,474.23,4850.2,1686.6,0.0000,7740.9,4449.7,4252.8,3658.0,0.0000,-620.83,-209.32,-125.83,-65.208,-203.74,-587.69,0.0000,-1105.4,-1695.4,-759.46,-1415.5
327.0000000000,192.88,2767.3,2908.9,2145.5,425.85,4410.6,1545.4,4.0752,6780.2,2555.0,3351.6,1976.2,0.0000,-9855.2,-8079.7,-2137.6,-3244.2,-4509.7,-18165.,-255.21,-21591.,-6486.1,-4596.7,-3226.4,94.885,3380.2,3082.2,2250.7,474.07,4850.2,1686.6,0.0000,7740.9,4449.7,4252.8,3658.0,0.0000,-620.27,-209.07,-125.80,-65.173,-203.84,-587.69,0.0000,-1105.3,-1694.9,-759.47,-1415.0
328.0000000000,192.84,2768.5,2909.5,2144.9,426.25,4410.4,1541.1,2.6899,6780.2,2555.6,3351.5,1976.7,0.0000,-9845.6,-8076.0,-2137.7,-3241.6,-4511.2,-18160.,-254.76,-21590.,-6486.4,-4596.9,-3225.5,105.75,3403.1,3108.1,2254.3,480.50,4852.4,1686.6,7.5268,7742.9,4451.7,4255.6,3660.9,0.0000,-623.13,-210.20,-126.13,-65.524,-203.94,-587.69,-0.34474,-1105.3,-1694.3,-759.49,-1414.7
329.0000000000,193.14,2777.9,2917.2,2144.8,427.85,4410.1,1482.1,2.6911,6780.3,2556.2,3351.5,1977.3,0.0000,-9837.1,-8072.9,-2137.8,-3239.0,-4512.6,-18155.,-254.32,-21590.,-6486.6,-4597.0,-3224.7,133.70,3443.5,3158.6,2261.4,495.34,4859.1,1686.6,11.617,7746.1,4454.4,4260.3,3666.0,0.0000,-627.19,-212.13,-126.57,-66.050,-204.07,-587.69,-0.53205,-1105.4,-1693.8,-759.52,-1414.6
330.0000000000,193.57,2788.3,2926.4,2145.7,429.56,4410.0,1461.6,2.6924,6747.3,2556.8,3351.4,1977.8,0.0000,-9829.5,-8070.4,-2138.0,-3236.6,-4513.8,-18151.,-253.86,-21589.,-6486.8,-4597.2,-3223.8,96.190,3426.7,3124.6,2256.5,480.16,4850.6,1686.6,0.0000,7740.9,4449.7,4252.8,3658.0,0.0000,-627.90,-211.52,-126.67,-66.045,-204.09,-587.69,0.0000,-1105.3,-1693.3,-759.49,-1413.5
331.0000000000,193.83,2792.8,2931.2,2146.5,430.48,4410.1,1418.9,2.6936,6673.4,2557.1,3351.4,1978.3,0.0000,-9822.3,-8067.9,-2138.1,-3234.2,-4514.8,-18146.,-253.40,-21588.,-6487.0,-4597.3,-3222.9,96.178,3426.3,3124.2,2256.4,480.10,4850.6,1686.6,0.0000,7740.9,4449.7,4252.8,3658.0,0.0000,-627.54,-211.36,-126.67,-66.029,-204.16,-587.69,0.0000,-1105.3,-1692.7,-759.50,-1413.0
332.0000000000,193.95,2793.6,2931.6,2146.7,430.65,4410.0,1418.9,2.6948,6591.7,2557.7,3351.4,1978.8,0.0000,-9815.1,-8065.4,-2138.2,-3231.8,-4515.7,-18142.,-252.94,-21587.,-6487.2,-4597.5,-3222.0,96.104,3423.7,3121.8,2256.1,479.76,4850.6,1686.6,0.0000,7740.9,4449.7,4252.8,3658.0,0.0000,-626.79,-211.07,-126.62,-65.971,-204.23,-587.69,0.0000,-1105.2,-1692.2,-759.51,-1412.6
333.0000000000,193.91,2792.7,2930.0,2146.7,430.43,4409.9,1377.7,2.6960,6577.1,2558.2,3351.5,1979.2,0.0000,-9807.7,-8062.9,-2138.3,-3229.3,-4516.3,-18137.,-252.48,-21587.,-6487.4,-4597.6,-3221.1,95.996,3419.8,3118.3,2255.6,479.25,4850.6,1686.6,0.0000,7740.9,4449.7,4252.8,3658.0,0.0000,-625.80,-210.70,-126.54,-65.888,-204.30,-587.69,0.0000,-1105.2,-1691.6,-759.52,-1412.1
334.0000000000,193.80,2790.8,2927.3,2146.1,430.00,4409.2,1355.5,2.6973,6576.9,2558.7,3351.5,1956.4,0.0000,-9800.2,-8060.2,-2138.3,-3226.8,-4516.8,-18133.,-252.02,-21586.,-6487.6,-4597.7,-3220.3,95.857,3414.8,3113.8,2251.5,478.54,4841.4,1686.6,0.0000,7735.3,4449.7,4252.8,3658.0,0.0000,-624.63,-210.27,-126.33,-65.784,-203.97,-587.69,0.0000,-1105.1,-1691.1,-759.52,-1411.6
335.0000000000,193.66,2788.4,2923.6,2144.7,429.36,4406.8,1355.5,2.6985,6576.2,2559.2,3351.5,1956.9,0.0000,-9792.5,-8057.5,-2138.2,-3224.4,-4517.0,-18128.,-251.56,-21585.,-6487.8,-4597.9,-3219.4,95.678,3408.5,3108.0,2246.8,477.64,4831.2,1686.6,0.0000,7729.1,4449.7,4252.8,3658.0,0.0000,-623.19,-209.75,-126.08,-65.652,-203.59,-587.69,0.0000,-1105.0,-1690.5,-759.53,-1411.1
336.0000000000,193.21,2784.9,2919.3,2142.4,428.62,4402.8,1355.5,2.6996,6575.1,2559.8,3351.5,1957.4,0.0000,-9784.7,-8054.6,-2138.1,-3221.9,-4516.9,-18124.,-251.10,-21584.,-6487.9,-4598.0,-3218.5,95.489,3401.7,3101.8,2242.0,476.69,4820.8,1686.6,0.0000,7722.9,4449.7,4252.8,3658.0,0.0000,-621.68,-209.20,-125.82,-65.513,-203.20,-587.69,0.0000,-1105.0,-1690.0,-759.54,-1410.6
337.0000000000,193.01,2780.9,2914.7,2139.0,427.74,4397.7,1355.5,2.6920,6573.4,2560.3,3351.4,1957.9,0.0000,-9776.5,-8051.6,-2137.8,-3219.3,-4516.5,-18119.,-250.65,-21583.,-6488.1,-4598.1,-3217.6,95.287,3394.5,3095.3,2237.0,475.68,4810.2,1686.6,0.0000,7716.5,4449.7,4252.8,3658.0,0.0000,-620.08,-208.62,-125.54,-65.365,-202.79,-587.69,0.0000,-1104.9,-1689.4,-759.55,-1410.1
338.0000000000,192.79,2776.3,2909.8,2135.0,426.85,4392.0,1355.6,2.6925,6571.1,2560.9,3351.4,1958.5,0.0000,-9768.2,-8048.6,-2137.5,-3216.8,-4515.8,-18115.,-250.20,-21582.,-6488.3,-4598.2,-3216.7,95.074,3387.0,3088.3,2231.9,474.62,4799.3,1686.6,0.0000,7709.9,4449.7,4252.8,3658.0,0.0000,-618.41,-208.02,-125.26,-65.209,-202.37,-587.69,0.0000,-1104.8,-1688.9,-759.55,-1409.6
339.0000000000,192.57,2771.8,2904.7,2130.7,425.95,4385.3,1355.6,2.6936,6567.6,2561.4,3351.4,1935.6,0.0000,-9759.6,-8045.4,-2137.0,-3214.3,-4514.8,-18110.,-249.74,-21580.,-6488.5,-4598.3,-3215.8,94.861,3379.4,3081.4,2226.8,473.55,4788.4,1686.6,0.0000,7703.3,4449.7,4252.8,3658.0,0.0000,-616.74,-207.41,-124.97,-65.053,-201.95,-587.69,0.0000,-1104.7,-1688.3,-759.56,-1409.1
340.0000000000,192.36,2767.8,2900.3,2126.5,425.26,4377.8,1355.5,1.7375,6563.2,2562.0,3351.4,1936.1,0.0000,-9751.0,-8042.3,-2136.6,-3211.8,-4513.7,-18106.,-249.29,-21579.,-6488.6,-4598.4,-3214.9,94.816,3377.8,3080.0,2224.9,473.31,4784.0,1686.6,0.0000,7700.6,4449.7,4252.8,3658.0,0.0000,-616.15,-207.17,-124.88,-65.011,-201.79,-587.69,0.0000,-1104.6,-1687.8,-759.57,-1408.6
341.0000000000,192.23,2764.6,2896.8,2122.8,424.72,4370.8,1355.5,0.85651,6558.8,2562.5,3351.4,1936.5,0.0000,-9742.5,-8039.1,-2136.0,-3209.2,-4512.3,-18101.,-248.84,-21577.,-6488.8,-4598.5,-3214.0,94.693,3373.4,3076.0,2221.2,472.68,4775.9,1686.6,0.0000,7695.7,4449.7,4252.8,3658.0,0.0000,-615.07,-206.76,-124.70,-64.917,-201.48,-587.69,0.0000,-1104.6,-1687.2,-759.57,-1408.1
342.0000000000,192.09,2761.2,2892.6,2119.5,424.25,4364.0,1303.0,0.85781,6554.4,2563.1,3351.4,1936.9,0.0000,-9733.9,-8036.0,-2135.5,-3206.7,-4510.9,-18097.,-248.40,-21577.,-6489.0,-4598.6,-3213.1,94.574,3369.2,3072.1,2217.7,472.08,4768.0,1686.6,0.0000,7691.0,4449.7,4252.8,3658.0,0.0000,-614.01,-206.36,-124.51,-64.826,-201.17,-587.69,0.0000,-1104.5,-1686.7,-759.58,-1407.6
343.0000000000,191.96,2757.5,2888.4,2116.2,423.68,4358.7,1292.1,0.85904,6549.9,2563.6,3351.3,1937.4,0.0000,-9725.2,-8032.8,-2134.9,-3204.2,-4509.2,-18092.,-247.95,-21579.,-6489.1,-4598.7,-3212.2,94.417,3363.6,3067.0,2213.5,471.29,4759.0,1686.6,0.0000,7685.5,4449.7,4252.8,3658.0,0.0000,-612.69,-205.88,-124.29,-64.708,-200.82,-587.69,0.0000,-1104.4,-1686.2,-759.59,-1407.1
344.0000000000,191.80,2753.9,2883.9,2112.8,423.04,4355.3,1292.1,0.86033,6545.4,2564.1,3351.2,1937.9,0.0000,-9716.5,-8029.7,-2134.3,-3201.7,-4507.4,-18088.,-247.50,-21580.,-6489.3,-4598.8,-3211.3,94.271,3358.4,3062.3,2209.5,470.55,4750.3,1686.6,0.0000,7680.2,4449.7,4252.8,3658.0,0.0000,-611.47,-205.42,-124.08,-64.598,-200.47,-587.69,0.0000,-1104.3,-1685.7,-759.59,-1406.6
345.0000000000,191.64,2749.8,2879.4,2109.2,422.37,4348.0,1245.4,0.86158,6541.4,2564.6,3351.1,1938.4,0.0000,-9707.7,-8026.4,-2133.6,-3199.2,-4505.4,-18083.,-247.05,-21581.,-6489.4,-4598.8,-3210.3,94.117,3352.9,3057.3,2205.4,469.77,4741.4,1686.6,0.0000,7674.8,4449.7,4252.8,3658.0,0.0000,-610.21,-204.94,-123.86,-64.483,-200.11,-587.69,0.0000,-1104.3,-1685.2,-759.60,-1406.1
346.0000000000,191.47,2745.7,2875.3,2105.5,421.68,4340.9,1165.9,0.86283,6537.3,2565.2,3351.1,1938.9,0.0000,-9698.8,-8023.2,-2132.9,-3196.7,-4503.2,-18079.,-246.61,-21581.,-6489.6,-4598.9,-3209.4,93.951,3347.0,3051.9,2201.1,468.94,4732.0,1686.6,0.0000,7669.2,4449.7,4252.8,3658.0,0.0000,-608.87,-204.43,-123.63,-64.359,-199.73,-587.69,0.0000,-1104.2,-1684.7,-759.60,-1405.6
347.0000000000,176.51,2741.7,2871.3,2101.7,420.99,4333.4,1165.9,0.86407,6533.1,2565.7,3351.1,1939.4,0.0000,-9689.9,-8019.9,-2132.2,-3194.2,-4500.9,-18075.,-246.16,-21580.,-6489.7,-4599.0,-3208.5,93.786,3341.1,3046.5,2196.8,468.10,4722.7,1686.6,0.0000,7663.5,4449.7,4252.8,3658.0,0.0000,-607.54,-203.93,-123.39,-64.236,-199.34,-587.69,0.0000,-1104.1,-1684.2,-759.61,-1405.1
348.0000000000,126.11,2737.4,2866.8,2098.0,420.27,4325.7,1165.9,0.86531,6528.6,2566.3,3351.1,1939.9,0.0000,-9681.0,-8016.5,-2131.4,-3191.7,-4498.3,-18070.,-245.72,-21579.,-6489.8,-4599.0,-3207.5,93.614,3334.9,3040.9,2192.4,467.24,4713.1,1686.6,0.0000,7657.8,4449.7,4252.8,3658.0,0.0000,-606.16,-203.41,-123.15,-64.108,-198.95,-587.69,0.0000,-1104.0,-1683.6,-759.61,-1404.6
349.0000000000,125.93,2732.7,2862.2,2094.1,419.54,4317.8,1165.9,0.86653,6523.9,2566.8,3351.1,1940.5,0.0000,-9672.0,-8013.1,-2130.5,-3189.2,-4495.6,-18066.,-245.27,-21578.,-6490.0,-4599.1,-3206.6,93.452,3329.2,3035.7,2188.1,466.42,4703.8,1686.6,0.0000,7652.1,4449.7,4252.8,3658.0,0.0000,-604.85,-202.91,-122.92,-63.987,-198.56,-587.69,0.0000,-1103.9,-1683.1,-759.62,-1404.1
350.0000000000,125.84,2728.2,2857.6,2090.1,418.82,4310.0,1165.9,0.86776,6519.2,2567.3,3351.1,1941.0,0.0000,-9662.9,-8009.7,-2129.7,-3186.7,-4492.8,-18061.,-244.83,-21577.,-6490.1,-4599.1,-3205.6,93.284,3323.2,3030.2,2183.7,465.58,4694.3,1686.6,0.0000,7646.4,4449.7,4252.8,3658.0,0.0000,-603.50,-202.39,-122.69,-63.862,-198.17,-587.69,0.0000,-1103.8,-1682.6,-759.62,-1403.6
351.0000000000,125.76,2723.4,2853.4,2086.0,418.08,4301.9,1144.9,0.86894,6514.3,2567.8,3351.1,1941.5,0.0000,-9653.8,-8006.3,-2128.8,-3184.1,-4489.7,-18057.,-244.39,-21575.,-6490.2,-4599.1,-3204.6,93.107,3316.9,3024.4,2179.2,464.68,4684.5,1686.6,0.0000,7640.5,4449.7,4252.8,3658.0,0.0000,-602.08,-201.86,-122.44,-63.730,-197.76,-587.69,0.0000,-1103.8,-1682.1,-759.63,-1403.1
352.0000000000,125.58,2718.3,2848.8,2082.0,417.31,4294.1,1102.5,0.87012,6509.0,2568.3,3351.1,1942.0,0.0000,-9644.6,-8003.0,-2127.8,-3181.6,-4486.6,-18053.,-243.95,-21574.,-6490.4,-4599.2,-3203.6,92.921,3310.3,3018.4,2174.5,463.75,4674.4,1686.6,0.0000,7634.4,4449.7,4252.8,3658.0,0.0000,-600.61,-201.30,-122.19,-63.592,-197.33,-587.69,0.0000,-1103.7,-1681.6,-759.63,-1402.6
353.0000000000,125.38,2713.4,2843.9,2077.8,416.51,4285.6,1102.5,0.87136,6503.8,2568.9,3351.0,1919.2,0.0000,-9635.2,-7999.5,-2126.8,-3179.1,-4483.2,-18048.,-243.51,-21572.,-6490.5,-4599.2,-3202.6,92.733,3303.6,3012.3,2169.8,462.81,4664.3,1686.6,0.0000,7628.2,4449.7,4252.8,3658.0,0.0000,-599.13,-200.74,-121.93,-63.453,-196.90,-587.69,0.0000,-1103.6,-1681.1,-759.64,-1402.1
354.0000000000,125.18,2708.6,2838.6,2073.5,415.69,4277.0,1102.5,0.87253,6498.6,2569.4,3351.0,1919.7,0.0000,-9625.8,-7996.1,-2125.8,-3176.6,-4479.8,-18044.,-243.07,-21571.,-6490.6,-4599.2,-3201.5,92.529,3296.3,3005.7,2164.8,461.79,4653.6,1686.6,0.0000,7621.8,4449.7,4252.8,3658.0,0.0000,-597.55,-200.15,-121.65,-63.304,-196.45,-587.69,0.0000,-1103.5,-1680.6,-759.64,-1401.5
355.0000000000,125.01,2705.9,2835.7,2069.4,415.34,4269.0,1081.0,0.87374,6493.5,2569.9,3351.0,1920.2,0.0000,-9616.5,-7992.8,-2124.8,-3174.1,-4476.2,-18039.,-242.64,-21569.,-6490.7,-4599.2,-3200.5,94.398,3304.9,3015.6,2167.1,464.43,4657.2,1686.6,0.25084,7623.8,4449.8,4253.3,3658.5,0.0000,-598.71,-200.53,-121.84,-63.456,-196.58,-587.69,-0.11489E-01,-1103.5,-1680.1,-759.65,-1401.1
356.0000000000,125.05,2707.0,2835.7,2066.7,415.41,4263.0,1039.1,0.87494,6488.9,2570.5,3351.0,1920.7,0.0000,-9607.6,-7989.7,-2123.8,-3171.6,-4472.6,-18035.,-242.21,-21567.,-6490.9,-4599.2,-3199.5,94.158,3304.4,3013.8,2165.0,463.25,4651.7,1686.6,0.0000,7620.5,4449.7,4252.8,3658.0,0.0000,-598.49,-200.36,-121.78,-63.443,-196.36,-587.69,0.0000,-1103.5,-1679.6,-759.65,-1400.5
357.0000000000,125.01,2706.2,2834.6,2064.7,415.43,4260.8,1039.1,0.87613,6484.6,2571.0,3351.1,1921.3,0.0000,-9598.9,-7986.6,-2122.9,-3169.2,-4468.9,-18031.,-241.78,-21566.,-6491.0,-4599.2,-3198.5,92.621,3299.6,3008.7,2162.2,462.16,4645.8,1686.6,0.0000,7617.0,4449.7,4252.8,3658.0,0.0000,-597.36,-199.91,-121.61,-63.339,-196.11,-587.69,0.0000,-1103.4,-1679.1,-759.66,-1400.0
358.0000000000,124.96,2703.1,2831.0,2062.7,415.03,4257.0,1039.1,0.87735,6480.2,2571.5,3351.1,1921.8,0.0000,-9590.1,-7983.2,-2121.9,-3166.7,-4465.3,-18026.,-241.35,-21564.,-6491.1,-4599.2,-3197.5,92.475,3294.4,3003.9,2160.8,461.47,4644.0,1686.6,0.0000,7616.0,4449.7,4252.8,3658.0,0.0000,-596.16,-199.45,-121.49,-63.230,-196.04,-587.69,0.0000,-1103.4,-1678.7,-759.66,-1399.4
359.0000000000,124.83,2699.6,2827.6,2060.9,414.42,4251.7,1039.1,0.87859,6476.4,2571.9,3351.1,1922.3,0.0000,-9581.2,-7979.9,-2121.0,-3164.3,-4461.5,-18022.,-240.91,-21562.,-6491.2,-4599.2,-3196.4,92.323,3289.0,2999.0,2159.5,460.75,4642.1,1686.6,0.0000,7614.9,4449.7,4252.8,3658.0,0.0000,-594.92,-198.97,-121.36,-63.116,-195.96,-587.69,0.0000,-1103.3,-1678.2,-759.66,-1398.9
360.0000000000,124.68,2696.7,2824.4,2059.2,413.90,4247.5,1039.1,0.87973,6473.8,2572.4,3351.1,1922.8,0.0000,-9572.4,-7976.6,-2120.1,-3161.8,-4457.8,-18018.,-240.48,-21561.,-6491.3,-4599.2,-3195.4,92.296,3288.0,2998.1,2159.0,460.62,4641.2,1686.6,0.0000,7614.3,4449.7,4252.8,3658.0,0.0000,-594.49,-198.77,-121.33,-63.089,-195.92,-587.69,0.0000,-1103.3,-1677.7,-759.67,-1398.4
361.0000000000,124.61,2696.2,2824.0,2057.7,413.83,4244.8,1039.0,0.88095,6471.7,2572.9,3351.0,1923.4,0.0000,-9563.8,-7973.4,-2119.2,-3159.4,-4454.0,-18013.,-240.05,-21559.,-6491.5,-4599.2,-3194.4,92.432,3295.3,3002.5,2160.7,461.25,4642.1,1686.6,1.1123,7615.2,4449.9,4252.8,3658.0,0.0000,-595.12,-198.92,-121.42,-63.172,-195.92,-587.69,-0.50943E-01,-1103.3,-1677.3,-759.67,-1397.8
362.0000000000,124.65,2698.3,2825.6,2057.0,414.16,4242.1,1039.0,0.88212,6407.8,2573.3,3351.0,1923.9,0.0000,-9555.6,-7970.5,-2118.4,-3157.0,-4450.2,-18009.,-239.63,-21557.,-6491.6,-4599.2,-3193.4,95.905,3301.8,3009.6,2161.9,462.02,4642.0,1686.6,1.5022,7615.4,4450.3,4253.1,3658.1,0.0000,-595.80,-199.15,-121.51,-63.263,-195.89,-587.69,-0.68801E-01,-1103.3,-1676.8,-759.68,-1397.3
363.0000000000,124.72,2699.6,2826.5,2056.9,414.37,4239.7,1039.0,0.88324,6398.4,2573.8,3350.9,1924.4,0.0000,-9547.6,-7967.7,-2117.6,-3154.7,-4446.4,-18005.,-239.20,-21555.,-6491.7,-4599.2,-3192.3,92.454,3293.6,3003.2,2158.8,461.34,4638.9,1686.6,0.0000,7612.8,4449.7,4252.8,3658.0,0.0000,-594.77,-198.70,-121.41,-63.171,-195.81,-587.69,0.0000,-1103.2,-1676.3,-759.68,-1396.7
364.0000000000,124.67,2698.2,2825.5,2056.4,414.22,4237.2,1039.0,0.88443,6396.7,2574.3,3350.9,1925.0,0.0000,-9539.6,-7964.9,-2116.7,-3152.3,-4442.6,-18000.,-238.77,-21553.,-6491.8,-4599.1,-3191.3,92.337,3289.5,2999.5,2157.6,460.78,4637.1,1686.6,0.0000,7611.8,4449.7,4252.8,3658.0,0.0000,-593.78,-198.32,-121.31,-63.083,-195.73,-587.69,0.0000,-1103.2,-1675.9,-759.68,-1396.2
365.0000000000,124.59,2695.9,2822.7,2055.4,413.78,4235.4,1038.9,0.88554,6395.3,2574.6,3350.9,1925.5,0.0000,-9531.6,-7962.0,-2115.9,-3149.9,-4438.7,-17996.,-238.34,-21551.,-6491.9,-4599.1,-3190.2,92.206,3284.8,2995.2,2156.3,460.16,4635.3,1686.6,0.0000,7610.7,4449.7,4252.8,3658.0,0.0000,-592.70,-197.90,-121.20,-62.985,-195.65,-587.69,0.0000,-1103.2,-1675.4,-759.68,-1395.6
366.0000000000,124.45,2692.9,2819.8,2054.4,413.24,4233.5,1038.9,0.88671,6393.9,2575.0,3350.9,1926.0,0.0000,-9523.4,-7959.1,-2115.1,-3147.6,-4434.8,-17992.,-237.92,-21550.,-6492.0,-4599.0,-3189.2,92.061,3279.6,2990.5,2155.0,459.47,4633.4,1686.6,0.0000,7609.6,4449.7,4252.8,3658.0,0.0000,-591.53,-197.46,-121.08,-62.877,-195.56,-587.69,0.0000,-1103.1,-1675.1,-759.69,-1395.1
367.0000000000,124.30,2689.3,2816.2,2053.3,412.66,4231.6,1038.9,0.88781,6392.6,2575.4,3351.0,1926.6,0.0000,-9515.2,-7956.1,-2114.3,-3145.2,-4430.8,-17987.,-237.49,-21548.,-6492.0,-4599.0,-3188.1,91.906,3274.1,2985.4,2153.5,458.73,4631.5,1686.6,0.0000,7608.5,4449.7,4252.8,3658.0,0.0000,-590.29,-196.99,-120.95,-62.762,-195.48,-587.69,0.0000,-1103.1,-1674.7,-759.69,-1394.5
368.0000000000,124.14,2685.8,2813.1,2052.1,412.05,4233.7,1038.9,0.88898,6391.2,2575.7,3350.9,1927.2,0.0000,-9506.8,-7953.1,-2113.5,-3142.8,-4426.9,-17983.,-237.06,-21546.,-6492.1,-4598.9,-3187.1,91.761,3268.9,2980.7,2152.2,458.04,4629.6,1686.6,0.0000,7607.4,4449.7,4252.8,3658.0,0.0000,-589.11,-196.54,-120.83,-62.654,-195.39,-587.69,0.0000,-1103.1,-1674.3,-759.69,-1393.9
369.0000000000,123.97,2682.1,2809.1,2051.1,411.34,4233.2,1038.8,0.89011,6389.9,2576.0,3350.9,1927.7,0.0000,-9498.4,-7950.1,-2112.6,-3140.4,-4422.8,-17979.,-236.64,-21544.,-6492.2,-4598.9,-3186.0,91.607,3263.4,2975.7,2150.8,457.31,4627.7,1686.6,0.0000,7606.2,4449.7,4252.8,3658.0,0.0000,-587.88,-196.08,-120.70,-62.540,-195.31,-587.69,0.0000,-1103.1,-1674.0,-759.69,-1393.4
370.0000000000,123.80,2678.1,2805.6,2049.9,410.70,4231.0,1038.8,0.89123,6388.5,2576.4,3350.9,1928.3,0.0000,-9489.9,-7947.0,-2111.8,-3138.0,-4418.8,-17974.,-236.22,-21542.,-6492.3,-4598.8,-3185.0,91.437,3257.4,2970.2,2149.3,456.51,4625.7,1686.6,0.0000,7605.0,4449.7,4252.8,3658.0,0.0000,-586.55,-195.58,-120.56,-62.414,-195.21,-587.69,0.0000,-1103.0,-1673.6,-759.70,-1392.8
371.0000000000,123.63,2674.2,2801.9,2048.6,410.09,4228.9,1038.8,0.89234,6387.0,2576.7,3350.9,1928.9,0.0000,-9481.3,-7943.9,-2111.0,-3135.6,-4414.7,-17970.,-235.79,-21540.,-6492.4,-4598.7,-3183.9,91.309,3252.8,2966.1,2148.1,455.90,4624.0,1686.6,0.0000,7604.0,4449.7,4252.8,3658.0,0.0000,-585.49,-195.17,-120.45,-62.318,-195.13,-587.69,0.0000,-1103.0,-1673.2,-759.70,-1392.3
372.0000000000,123.48,2670.8,2798.2,2047.3,409.55,4227.0,985.80,0.89346,6385.7,2577.1,3350.9,1929.4,0.0000,-9472.7,-7940.8,-2110.1,-3133.2,-4410.6,-17966.,-235.37,-21538.,-6492.4,-4598.6,-3182.9,91.201,3249.0,2962.5,2147.0,455.39,4622.3,1686.6,0.0000,7603.0,4449.7,4252.8,3658.0,0.0000,-584.55,-194.80,-120.36,-62.235,-195.06,-587.69,0.0000,-1103.0,-1672.9,-759.70,-1391.7
373.0000000000,123.34,2667.6,2794.8,2046.0,409.05,4225.0,975.05,0.89457,6384.5,2577.5,3350.9,1930.0,0.0000,-9464.1,-7937.7,-2109.3,-3130.8,-4406.5,-17962.,-234.95,-21536.,-6492.5,-4598.5,-3181.8,91.071,3244.4,2958.3,2145.7,454.77,4620.6,1686.6,0.0000,7602.0,4449.7,4252.8,3658.0,0.0000,-583.47,-194.38,-120.25,-62.137,-194.97,-587.69,0.0000,-1102.9,-1672.5,-759.70,-1391.2
374.0000000000,123.20,2663.9,2791.0,2044.8,408.51,4222.9,975.04,0.89567,6383.2,2577.8,3350.9,1930.5,0.0000,-9455.5,-7934.6,-2108.4,-3128.4,-4402.3,-17957.,-234.53,-21534.,-6492.6,-4598.5,-3180.8,90.901,3238.3,2952.8,2144.2,453.96,4618.6,1686.6,0.0000,7600.8,4449.7,4252.8,3658.0,0.0000,-582.14,-193.88,-120.11,-62.012,-194.88,-587.69,0.0000,-1102.9,-1672.1,-759.70,-1390.6
375.0000000000,123.03,2659.7,2786.5,2043.5,407.87,4220.9,975.03,0.89673,6382.0,2578.2,3350.9,1931.0,0.0000,-9446.8,-7931.4,-2107.5,-3126.1,-4398.1,-17953.,-234.11,-21532.,-6492.6,-4598.4,-3179.7,90.721,3231.9,2946.9,2142.6,453.11,4616.5,1686.6,0.0000,7599.6,4449.7,4252.8,3658.0,0.0000,-580.74,-193.36,-119.97,-61.879,-194.78,-587.69,0.0000,-1102.9,-1671.8,-759.71,-1390.1
376.0000000000,122.96,2655.0,2781.4,2042.2,407.15,4219.0,975.03,0.89783,6380.9,2578.5,3350.9,1931.6,0.0000,-9438.0,-7928.1,-2106.7,-3123.7,-4393.9,-17949.,-233.69,-21530.,-6492.7,-4598.3,-3178.7,90.532,3225.2,2940.8,2141.0,452.21,4614.4,1686.6,0.0000,7598.3,4449.7,4252.8,3658.0,0.0000,-579.29,-192.82,-119.81,-61.741,-194.68,-587.69,0.0000,-1102.8,-1671.4,-759.71,-1389.5
377.0000000000,122.64,2650.2,2775.9,2040.9,406.40,4217.0,975.00,0.89896,6379.7,2578.9,3350.8,1932.1,0.0000,-9429.1,-7924.7,-2105.8,-3121.3,-4389.7,-17944.,-233.28,-21528.,-6492.7,-4598.2,-3177.6,90.338,3218.2,2934.5,2139.3,451.29,4612.2,1686.6,0.0000,7597.1,4449.7,4252.8,3658.0,0.0000,-577.80,-192.26,-119.65,-61.599,-194.58,-587.69,0.0000,-1102.8,-1671.0,-759.71,-1389.0
378.0000000000,122.36,2645.1,2770.4,2039.5,405.62,4215.0,974.97,0.90004,6378.5,2579.3,3350.8,1932.7,0.0000,-9420.0,-7921.3,-2104.9,-3118.9,-4385.4,-17940.,-232.86,-21526.,-6492.8,-4598.0,-3176.5,90.141,3211.2,2928.1,2137.6,450.36,4610.0,1686.6,0.0000,7595.8,4449.7,4252.8,3658.0,0.0000,-576.29,-191.70,-119.50,-61.455,-194.48,-587.69,0.0000,-1102.8,-1670.7,-759.71,-1388.4
379.0000000000,122.17,2640.1,2764.9,2038.0,404.86,4213.2,974.96,0.90112,6377.4,2579.6,3350.8,1933.2,0.0000,-9410.9,-7917.8,-2104.0,-3116.5,-4381.1,-17936.,-232.44,-21524.,-6492.8,-4597.9,-3175.5,89.972,3205.2,2922.6,2136.4,449.56,4608.7,1686.6,0.0000,7595.0,4449.7,4252.8,3658.0,0.0000,-574.96,-191.19,-119.37,-61.330,-194.41,-587.69,0.0000,-1102.7,-1670.3,-759.71,-1387.9
380.0000000000,121.82,2635.4,2760.2,2036.7,404.14,4211.3,974.91,0.90220,6376.2,2580.0,3350.9,1933.7,0.0000,-9401.7,-7914.4,-2103.1,-3114.1,-4376.8,-17932.,-232.03,-21522.,-6492.9,-4597.8,-3174.4,89.801,3199.1,2917.0,2135.5,448.76,4608.4,1686.6,0.0000,7594.8,4449.7,4252.8,3658.0,0.0000,-573.61,-190.69,-119.25,-61.204,-194.39,-587.69,0.0000,-1102.7,-1669.9,-759.71,-1387.4
381.0000000000,121.53,2630.7,2755.3,2035.6,403.47,4209.9,974.91,0.90327,6375.2,2580.3,3350.9,1934.3,0.0000,-9392.5,-7910.9,-2102.1,-3111.7,-4372.5,-17927.,-231.62,-21521.,-6492.9,-4597.7,-3173.4,89.641,3193.4,2911.9,2134.7,448.01,4608.1,1686.6,0.0000,7594.7,4449.7,4252.8,3658.0,0.0000,-572.34,-190.20,-119.14,-61.085,-194.37,-587.69,0.0000,-1102.6,-1669.6,-759.71,-1386.8
382.0000000000,121.35,2626.2,2750.5,2034.6,402.79,4208.8,974.87,0.90433,6374.2,2580.7,3350.8,1934.8,0.0000,-9383.2,-7907.5,-2101.2,-3109.3,-4368.2,-17923.,-231.20,-21519.,-6492.9,-4597.5,-3172.3,89.464,3187.1,2906.1,2133.8,447.19,4607.8,1686.6,0.0000,7594.5,4449.7,4252.8,3658.0,0.0000,-570.96,-189.68,-119.02,-60.956,-194.34,-587.69,0.0000,-1102.6,-1669.2,-759.71,-1386.3
383.0000000000,121.17,2621.5,2745.7,2033.7,402.12,4207.7,974.86,0.90540,6373.3,2581.1,3350.8,1935.4,0.0000,-9373.9,-7904.0,-2100.3,-3106.9,-4363.9,-17919.,-230.79,-21516.,-6492.9,-4597.4,-3171.2,89.297,3181.2,2900.7,2133.0,446.40,4607.4,1686.6,0.0000,7594.4,4449.7,4252.8,3658.0,0.0000,-569.64,-189.18,-118.90,-60.832,-194.32,-587.69,0.0000,-1102.5,-1668.8,-759.71,-1385.7
384.0000000000,120.99,2616.7,2740.8,2032.8,401.43,4206.7,974.85,0.90642,6372.6,2581.4,3350.8,1935.9,0.0000,-9364.6,-7900.5,-2099.5,-3104.5,-4359.6,-17915.,-230.38,-21514.,-6493.0,-4597.3,-3170.2,89.118,3174.8,2894.9,2132.0,445.57,4607.1,1686.6,0.0000,7594.2,4449.7,4252.8,3658.0,0.0000,-568.25,-188.65,-118.78,-60.700,-194.29,-587.69,0.0000,-1102.5,-1668.5,-759.71,-1385.2
385.0000000000,120.80,2611.9,2735.6,2031.9,400.73,4205.9,974.85,0.90751,6372.1,2581.8,3350.8,1936.5,0.0000,-9355.2,-7897.0,-2098.6,-3102.1,-4355.3,-17910.,-229.97,-21512.,-6493.0,-4597.1,-3169.1,88.930,3168.1,2888.8,2131.1,444.69,4606.8,1686.6,0.0000,7594.0,4449.7,4252.8,3658.0,0.0000,-566.80,-188.11,-118.65,-60.563,-194.26,-587.69,0.0000,-1102.4,-1668.1,-759.71,-1384.7
386.0000000000,120.60,2607.0,2730.1,2031.0,399.99,4205.3,974.85,0.90857,6371.8,2582.2,3350.8,1937.0,0.0000,-9345.7,-7893.5,-2097.7,-3099.7,-4351.0,-17906.,-229.56,-21510.,-6493.0,-4596.9,-3168.1,88.735,3161.1,2882.4,2130.1,443.78,4606.4,1686.6,0.0000,7593.9,4449.7,4252.8,3658.0,0.0000,-565.30,-187.55,-118.52,-60.420,-194.24,-587.69,0.0000,-1102.4,-1667.7,-759.71,-1384.1
387.0000000000,120.40,2602.0,2724.7,2030.1,399.27,4204.5,974.84,0.90961,6371.5,2582.5,3350.8,1937.6,0.0000,-9336.2,-7889.9,-2096.8,-3097.3,-4346.7,-17902.,-229.15,-21508.,-6493.0,-4596.8,-3167.0,88.570,3155.3,2877.1,2129.3,443.01,4606.1,1686.6,0.0000,7593.7,4449.7,4252.8,3658.0,0.0000,-563.99,-187.05,-118.40,-60.298,-194.21,-587.69,0.0000,-1102.3,-1667.4,-759.71,-1383.6
388.0000000000,120.21,2597.3,2719.3,2029.2,398.57,4204.0,974.84,0.91062,6371.3,2582.9,3350.8,1938.1,0.0000,-9326.6,-7886.4,-2095.9,-3094.9,-4342.4,-17898.,-228.74,-21506.,-6493.0,-4596.6,-3165.9,88.396,3149.1,2871.4,2128.4,442.19,4605.8,1686.6,0.0000,7593.6,4449.7,4252.8,3658.0,0.0000,-562.63,-186.53,-118.28,-60.170,-194.19,-587.69,0.0000,-1102.2,-1667.0,-759.71,-1383.1
389.0000000000,120.03,2593.0,2714.5,2028.4,397.98,4203.3,974.82,0.91166,6371.0,2583.2,3350.8,1938.5,0.0000,-9317.1,-7882.8,-2095.0,-3092.5,-4338.1,-17893.,-228.34,-21504.,-6493.0,-4596.4,-3164.9,88.304,3145.8,2868.4,2127.9,441.76,4605.6,1686.6,0.0000,7593.4,4449.7,4252.8,3658.0,0.0000,-561.79,-186.19,-118.22,-60.098,-194.16,-587.69,0.0000,-1102.2,-1666.7,-759.72,-1382.6
390.0000000000,119.89,2589.5,2710.5,2027.6,397.48,4202.8,974.79,0.91269,6370.8,2583.6,3350.7,1939.0,0.0000,-9307.6,-7879.3,-2094.1,-3090.1,-4333.7,-17889.,-227.93,-21502.,-6493.0,-4596.3,-3163.8,88.178,3141.3,2864.3,2127.3,441.17,4605.3,1686.6,0.0000,7593.3,4449.7,4252.8,3658.0,0.0000,-560.73,-185.77,-118.13,-60.003,-194.14,-587.69,0.0000,-1102.1,-1666.3,-759.72,-1382.0
391.0000000000,119.74,2585.8,2706.2,2026.9,396.96,4202.4,974.79,0.91376,6370.5,2584.0,3350.7,1939.5,0.0000,-9298.1,-7875.9,-2093.2,-3087.7,-4329.4,-17885.,-227.53,-21500.,-6493.0,-4596.1,-3162.7,88.012,3135.4,2858.9,2126.4,440.39,4605.0,1686.6,0.0000,7593.1,4449.7,4252.8,3658.0,0.0000,-559.42,-185.28,-118.02,-59.881,-194.11,-587.69,0.0000,-1102.1,-1665.9,-759.73,-1381.5
392.0000000000,119.58,2581.3,2701.3,2026.2,396.33,4201.9,974.79,0.91478,6370.3,2584.3,3350.6,1940.1,0.0000,-9288.6,-7872.3,-2092.3,-3085.3,-4325.0,-17881.,-227.12,-21498.,-6493.0,-4595.9,-3161.7,87.816,3128.4,2852.6,2125.4,439.48,4604.6,1686.6,0.0000,7592.9,4449.7,4252.8,3658.0,0.0000,-557.93,-184.72,-117.88,-59.738,-194.08,-587.69,0.0000,-1102.0,-1665.6,-759.73,-1381.0
393.0000000000,119.40,2576.7,2696.5,2025.5,395.68,4201.5,974.76,0.91577,6370.2,2584.7,3350.6,1940.6,0.0000,-9279.0,-7868.8,-2091.4,-3083.0,-4320.7,-17877.,-226.72,-21496.,-6493.0,-4595.7,-3160.6,87.685,3123.7,2848.3,2124.7,438.87,4604.3,1686.6,0.0000,7592.8,4449.7,4252.8,3658.0,0.0000,-556.84,-184.29,-117.79,-59.640,-194.05,-587.69,0.0000,-1102.0,-1665.2,-759.74,-1380.5
394.0000000000,119.24,2572.8,2692.2,2024.7,395.12,4201.1,974.74,0.91682,6370.1,2585.0,3350.6,1941.1,0.0000,-9269.5,-7865.3,-2090.5,-3080.6,-4316.3,-17872.,-226.31,-21494.,-6493.0,-4595.5,-3159.5,87.578,3119.9,2844.9,2124.2,438.37,4604.1,1686.6,0.0000,7592.7,4449.7,4252.8,3658.0,0.0000,-555.91,-183.92,-117.72,-59.558,-194.03,-587.69,0.0000,-1101.9,-1664.9,-759.74,-1380.0
395.0000000000,119.09,2569.4,2687.7,2024.0,394.63,4200.7,974.70,0.91783,6369.9,2585.4,3350.6,1941.6,0.0000,-9260.1,-7861.8,-2089.7,-3078.2,-4312.0,-17868.,-225.91,-21492.,-6493.0,-4595.3,-3158.5,87.456,3115.6,2840.9,2123.5,437.79,4603.8,1686.6,0.0000,7592.5,4449.7,4252.8,3658.0,0.0000,-554.88,-183.52,-117.63,-59.465,-194.00,-587.69,0.0000,-1101.8,-1664.5,-759.75,-1379.4
396.0000000000,118.95,2565.7,2682.8,2023.3,394.10,4200.3,974.69,0.93172,6369.7,2585.7,3350.6,1942.2,0.0000,-9250.6,-7858.4,-2088.8,-3075.9,-4307.6,-17864.,-225.51,-21489.,-6493.0,-4595.1,-3157.4,87.280,3109.3,2835.2,2122.6,436.97,4603.4,1686.6,0.0000,7592.3,4449.7,4252.8,3658.0,0.0000,-553.52,-183.00,-117.51,-59.337,-193.97,-587.69,0.0000,-1101.8,-1664.2,-759.75,-1378.9
397.0000000000,118.78,2561.1,2677.7,2022.6,393.42,4200.0,974.68,0.93937,6369.6,2586.1,3350.6,1942.7,0.0000,-9241.1,-7854.9,-2087.9,-3073.5,-4303.2,-17860.,-225.11,-21487.,-6492.9,-4594.8,-3156.3,87.077,3102.1,2828.6,2121.7,436.02,4603.3,1686.6,0.0000,7592.3,4449.7,4252.8,3658.0,0.0000,-551.98,-182.43,-117.38,-59.190,-193.95,-587.69,0.0000,-1101.7,-1663.8,-759.76,-1378.4
398.0000000000,118.59,2556.1,2671.5,2021.9,392.67,4199.6,974.68,0.94039,6369.4,2586.5,3350.5,1943.2,0.0000,-9231.5,-7851.4,-2087.0,-3071.2,-4298.9,-17856.,-224.71,-21485.,-6492.9,-4594.6,-3155.3,86.876,3094.9,2822.0,2120.8,435.08,4603.2,1686.6,0.0000,7592.3,4449.7,4252.8,3658.0,0.0000,-550.46,-181.86,-117.24,-59.044,-193.93,-587.69,0.0000,-1101.7,-1663.5,-759.76,-1377.9
399.0000000000,118.38,2551.3,2665.8,2021.1,391.95,4199.3,974.66,0.94140,6369.3,2586.8,3350.4,1943.7,0.0000,-9221.8,-7847.8,-2086.1,-3068.8,-4294.5,-17851.,-224.31,-21483.,-6492.9,-4594.4,-3154.2,86.735,3089.9,2817.5,2120.2,434.43,4603.2,1686.6,0.0000,7592.3,4449.7,4252.8,3658.0,0.0000,-549.31,-181.41,-117.15,-58.939,-193.91,-587.69,0.0000,-1101.6,-1663.1,-759.76,-1377.4
400.0000000000,118.21,2547.1,2660.9,2020.4,391.32,4199.0,974.65,0.94241,6369.1,2587.2,3350.4,1944.2,0.0000,-9212.2,-7844.3,-2085.2,-3066.5,-4290.1,-17847.,-223.92,-21481.,-6492.9,-4594.1,-3153.1,86.585,3084.5,2812.6,2119.5,433.73,4603.1,1686.6,0.0000,7592.3,4449.7,4252.8,3658.0,0.0000,-548.11,-180.95,-117.05,-58.827,-193.89,-587.69,0.0000,-1101.6,-1662.8,-759.77,-1376.9
401.0000000000,118.03,2542.8,2656.3,2019.7,390.71,4198.7,974.65,0.94341,6369.0,2587.5,3350.4,1944.7,0.0000,-9202.6,-7840.7,-2084.3,-3064.1,-4285.8,-17843.,-223.52,-21479.,-6492.8,-4593.9,-3152.0,86.409,3078.3,2806.9,2118.7,432.90,4603.0,1686.6,0.0000,7592.3,4449.7,4252.8,3658.0,0.0000,-546.74,-180.44,-116.93,-58.698,-193.87,-587.69,0.0000,-1101.5,-1662.4,-759.77,-1376.4
402.0000000000,117.86,2538.6,2651.9,2019.1,390.12,4198.5,974.64,0.94441,6368.9,2587.9,3350.4,1945.2,0.0000,-9192.9,-7837.3,-2083.4,-3061.8,-4281.4,-17839.,-223.12,-21476.,-6492.8,-4593.7,-3151.0,86.292,3074.1,2803.1,2118.2,432.36,4603.0,1686.6,0.0000,7592.3,4449.7,4252.8,3658.0,0.0000,-545.76,-180.04,-116.85,-58.610,-193.85,-587.69,0.0000,-1101.5,-1662.1,-759.78,-1375.9
403.0000000000,117.71,2535.0,2647.9,2018.5,389.61,4198.2,974.64,0.94541,6368.8,2588.2,3350.4,1945.7,0.0000,-9183.3,-7833.9,-2082.5,-3059.4,-4277.0,-17835.,-222.73,-21474.,-6492.7,-4593.4,-3149.9,86.184,3070.3,2799.6,2117.7,431.86,4602.9,1686.6,0.0000,7592.3,4449.7,4252.8,3658.0,0.0000,-544.82,-179.67,-116.78,-58.528,-193.84,-587.69,0.0000,-1101.4,-1661.7,-759.78,-1375.4
404.0000000000,117.57,2531.7,2644.1,2017.9,389.11,4198.0,974.64,0.94639,6368.7,2588.6,3350.4,1946.2,0.0000,-9173.8,-7830.5,-2081.6,-3057.1,-4272.7,-17831.,-222.33,-21472.,-6492.7,-4593.2,-3148.8,86.050,3065.5,2795.2,2117.1,431.23,4602.9,1686.6,0.0000,7592.2,4449.7,4252.8,3658.0,0.0000,-543.72,-179.25,-116.69,-58.428,-193.82,-587.69,0.0000,-1101.3,-1661.4,-759.78,-1374.9
405.0000000000,117.43,2527.7,2639.8,2017.3,388.54,4197.8,974.63,0.94739,6368.7,2588.9,3350.4,1946.7,0.0000,-9164.3,-7827.1,-2080.7,-3054.8,-4268.3,-17827.,-221.94,-21470.,-6492.7,-4592.9,-3147.7,85.867,3059.0,2789.3,2116.3,430.38,4602.8,1686.6,0.0000,7592.2,4449.7,4252.8,3658.0,0.0000,-542.32,-178.72,-116.57,-58.295,-193.80,-587.69,0.0000,-1101.3,-1661.0,-759.79,-1374.4
406.0000000000,117.25,2523.0,2634.5,2016.7,387.85,4197.6,974.63,0.94836,6369.0,2589.3,3350.4,1947.2,0.0000,-9154.7,-7823.6,-2079.8,-3052.4,-4263.9,-17823.,-221.55,-21467.,-6492.6,-4592.6,-3146.7,85.666,3051.8,2782.7,2115.3,429.44,4602.7,1686.6,0.0000,7592.2,4449.7,4252.8,3658.0,0.0000,-540.80,-178.15,-116.44,-58.149,-193.78,-587.69,0.0000,-1101.2,-1660.7,-759.79,-1373.9
407.0000000000,117.01,2518.3,2629.5,2016.1,387.16,4197.3,974.63,0.94935,6369.0,2589.6,3350.4,1947.7,0.0000,-9145.1,-7820.1,-2078.9,-3050.1,-4259.6,-17818.,-221.15,-21465.,-6492.5,-4592.4,-3145.6,85.533,3047.1,2778.4,2114.7,428.82,4602.6,1686.6,0.0000,7592.2,4449.7,4252.8,3658.0,0.0000,-539.71,-177.73,-116.35,-58.050,-193.75,-587.69,0.0000,-1101.2,-1660.3,-759.79,-1373.4
408.0000000000,116.61,2514.3,2625.2,2015.4,386.58,4197.2,974.63,0.95032,6369.0,2590.0,3350.4,1948.1,0.0000,-9135.5,-7816.6,-2078.0,-3047.8,-4255.2,-17814.,-220.76,-21463.,-6492.5,-4592.1,-3144.5,85.419,3043.0,2774.7,2114.2,428.28,4602.6,1686.6,0.0000,7592.2,4449.7,4252.8,3658.0,0.0000,-538.75,-177.35,-116.27,-57.964,-193.73,-587.69,0.0000,-1101.1,-1660.0,-759.79,-1372.9
409.0000000000,116.45,2510.5,2620.8,2014.8,386.03,4197.0,974.62,0.95130,6369.1,2590.4,3350.4,1948.6,0.0000,-9126.0,-7813.2,-2077.1,-3045.5,-4250.8,-17810.,-220.37,-21461.,-6492.4,-4591.8,-3143.4,85.252,3037.1,2769.3,2113.5,427.50,4602.5,1686.6,0.0000,7592.2,4449.7,4252.8,3658.0,0.0000,-537.45,-176.85,-116.16,-57.841,-193.71,-587.69,0.0000,-1101.1,-1659.6,-759.80,-1372.5
410.0000000000,116.28,2506.0,2616.0,2014.3,385.39,4196.9,974.62,0.95227,6369.1,2590.7,3350.4,1949.1,0.0000,-9116.4,-7809.7,-2076.2,-3043.2,-4246.5,-17806.,-219.98,-21458.,-6492.4,-4591.5,-3142.3,85.057,3030.1,2763.0,2112.6,426.59,4602.4,1686.6,0.0000,7592.2,4449.7,4252.8,3658.0,0.0000,-535.97,-176.30,-116.03,-57.700,-193.69,-587.69,0.0000,-1101.0,-1659.3,-759.80,-1372.0
411.0000000000,116.12,2500.9,2610.6,2013.6,384.64,4196.8,974.62,0.95323,6369.1,2591.1,3350.4,1949.6,0.0000,-9106.7,-7806.2,-2075.3,-3040.9,-4242.1,-17802.,-219.60,-21456.,-6492.3,-4591.2,-3141.3,84.843,3022.5,2756.0,2111.6,425.60,4602.3,1686.6,0.0000,7592.2,4449.7,4252.8,3658.0,0.0000,-534.38,-175.72,-115.89,-57.546,-193.67,-587.69,0.0000,-1101.0,-1658.9,-759.80,-1371.5
412.0000000000,115.92,2495.3,2605.2,2012.8,383.82,4196.7,974.62,0.95419,6369.2,2591.4,3350.4,1950.1,0.0000,-9096.9,-7802.7,-2074.3,-3038.5,-4237.8,-17798.,-219.21,-21454.,-6492.2,-4590.9,-3140.2,84.628,3014.8,2749.0,2110.7,424.59,4602.2,1686.6,0.0000,7592.2,4449.7,4252.8,3658.0,0.0000,-532.78,-175.12,-115.74,-57.391,-193.65,-587.69,0.0000,-1100.9,-1658.6,-759.80,-1371.0
413.0000000000,115.70,2489.6,2599.4,2012.0,382.97,4196.6,974.61,0.95514,6369.2,2591.8,3350.3,1949.6,0.0000,-9087.1,-7799.1,-2073.4,-3036.2,-4233.4,-17794.,-218.82,-21451.,-6492.2,-4590.7,-3139.1,84.406,3006.9,2741.8,2109.7,423.56,4602.2,1686.6,0.0000,7592.2,4449.7,4252.8,3658.0,0.0000,-531.13,-174.52,-115.59,-57.232,-193.63,-587.69,0.0000,-1100.9,-1658.2,-759.80,-1370.5
414.0000000000,115.47,2483.8,2593.4,2011.2,382.10,4196.4,974.61,0.95606,6369.2,2592.1,3350.2,1951.1,0.0000,-9077.1,-7795.4,-2072.5,-3033.9,-4229.1,-17790.,-218.44,-21449.,-6492.1,-4590.4,-3138.0,84.182,2999.0,2734.5,2108.7,422.51,4602.1,1686.6,0.0000,7592.2,4449.7,4252.8,3658.0,0.0000,-529.47,-173.90,-115.44,-57.070,-193.61,-587.69,0.0000,-1100.8,-1657.9,-759.81,-1370.1
415.0000000000,115.23,2477.7,2587.3,2010.4,381.21,4196.3,974.60,0.95701,6369.3,2592.5,3350.2,1951.5,0.0000,-9067.1,-7791.7,-2071.6,-3031.5,-4224.7,-17786.,-218.05,-21447.,-6492.0,-4590.0,-3136.9,83.950,2990.7,2727.0,2107.6,421.43,4602.0,1686.6,0.0000,7592.2,4449.7,4252.8,3658.0,0.0000,-527.76,-173.27,-115.29,-56.904,-193.59,-587.69,0.0000,-1100.7,-1657.6,-759.81,-1369.6
416.0000000000,114.99,2471.5,2580.8,2009.7,380.30,4196.2,974.56,0.95799,6369.3,2592.8,3350.2,1952.0,0.0000,-9057.0,-7788.0,-2070.6,-3029.2,-4220.4,-17782.,-217.67,-21444.,-6492.0,-4589.7,-3135.9,83.710,2982.1,2719.2,2106.6,420.31,4601.9,1686.6,0.0000,7592.2,4449.7,4252.8,3658.0,0.0000,-526.00,-172.63,-115.13,-56.731,-193.57,-587.69,0.0000,-1100.7,-1657.2,-759.81,-1369.1
417.0000000000,114.75,2465.4,2574.3,2008.8,379.41,4196.0,974.56,0.95890,6369.4,2593.1,3350.2,1929.2,0.0000,-9046.8,-7784.3,-2069.7,-3026.9,-4216.0,-17778.,-217.28,-21442.,-6491.9,-4589.4,-3134.8,83.512,2975.1,2712.8,2105.7,419.38,4601.9,1686.6,0.0000,7592.2,4449.7,4252.8,3658.0,0.0000,-524.50,-172.07,-115.00,-56.588,-193.55,-587.69,0.0000,-1100.6,-1656.9,-759.81,-1368.6
418.0000000000,114.52,2459.8,2568.3,2007.9,378.59,4195.9,974.56,0.95987,6369.4,2593.5,3350.2,1929.6,0.0000,-9036.5,-7780.5,-2068.8,-3024.5,-4211.7,-17774.,-216.90,-21440.,-6491.8,-4589.1,-3133.7,83.325,2968.4,2706.7,2104.8,418.51,4601.8,1686.6,0.0000,7592.2,4449.7,4252.8,3658.0,0.0000,-523.08,-171.53,-114.87,-56.452,-193.52,-587.69,0.0000,-1100.6,-1656.5,-759.81,-1368.2
419.0000000000,114.30,2454.2,2562.3,2007.1,377.77,4195.8,974.55,0.96080,6369.5,2593.8,3350.2,1930.1,0.0000,-9026.2,-7776.7,-2067.8,-3022.2,-4207.3,-17770.,-216.52,-21437.,-6491.7,-4588.8,-3132.6,83.093,2960.2,2699.2,2103.8,417.43,4601.7,1686.6,0.0000,7592.1,4449.7,4252.8,3658.0,0.0000,-521.37,-170.90,-114.72,-56.286,-193.50,-587.69,0.0000,-1100.5,-1656.2,-759.81,-1367.7
420.0000000000,114.07,2448.0,2555.9,2006.3,376.86,4195.5,974.55,0.96172,6369.5,2594.1,3350.2,1930.6,0.0000,-9015.9,-7772.9,-2066.9,-3019.8,-4203.0,-17766.,-216.14,-21435.,-6491.7,-4588.5,-3131.5,82.845,2951.3,2691.1,2102.7,416.27,4601.6,1686.6,0.0000,7592.1,4449.7,4252.8,3658.0,0.0000,-519.56,-170.24,-114.55,-56.108,-193.48,-587.69,0.0000,-1100.5,-1655.9,-759.81,-1367.2
421.0000000000,113.84,2441.2,2549.1,2005.5,375.85,4195.4,974.51,0.97725,6369.6,2594.4,3350.2,1931.1,0.0000,-9005.5,-7769.1,-2065.9,-3017.5,-4198.6,-17762.,-215.76,-21433.,-6491.6,-4588.1,-3130.5,82.608,2942.9,2683.4,2101.6,415.17,4601.6,1686.6,0.0000,7592.1,4449.7,4252.8,3658.0,0.0000,-517.82,-169.60,-114.40,-55.938,-193.46,-587.69,0.0000,-1100.4,-1655.6,-759.81,-1366.7
422.0000000000,113.72,2437.7,2545.4,2004.7,375.51,4195.3,974.50,0.97867,6369.7,2594.8,3350.2,1931.6,0.0000,-8995.2,-7765.3,-2065.0,-3015.2,-4194.3,-17758.,-215.38,-21430.,-6491.5,-4587.8,-3129.4,82.974,2954.3,2693.7,2103.2,416.74,4601.7,1686.6,0.0000,7592.1,4449.7,4252.8,3658.0,0.0000,-519.53,-170.09,-114.60,-56.142,-193.44,-587.69,0.0000,-1100.4,-1655.2,-759.81,-1366.2
423.0000000000,113.85,2439.3,2546.1,2004.1,375.75,4195.2,974.50,0.97960,6369.8,2595.1,3350.2,1932.1,0.0000,-8985.6,-7761.9,-2064.1,-3012.9,-4190.0,-17754.,-215.01,-21428.,-6491.4,-4587.5,-3128.3,82.959,2955.4,2694.8,2103.2,416.80,4601.7,1686.6,0.0000,7592.1,4449.7,4252.8,3658.0,0.0000,-519.52,-170.02,-114.63,-56.159,-193.41,-587.69,0.0000,-1100.3,-1654.9,-759.81,-1365.8
424.0000000000,113.81,2439.2,2545.8,2004.1,375.89,4195.2,974.48,0.98050,6369.8,2595.4,3350.1,1932.5,0.0000,-8976.2,-7758.6,-2063.2,-3010.7,-4185.6,-17750.,-214.63,-21425.,-6491.3,-4587.1,-3127.2,82.839,2951.1,2690.9,2102.7,416.24,4601.6,1686.6,0.0000,7592.1,4449.7,4252.8,3658.0,0.0000,-518.53,-169.64,-114.55,-56.070,-193.39,-587.69,0.0000,-1100.3,-1654.6,-759.81,-1365.3
425.0000000000,113.81,2436.3,2542.9,2003.9,375.65,4195.0,974.42,0.98142,6369.8,2595.8,3350.1,1933.0,0.0000,-8966.9,-7755.4,-2062.3,-3008.5,-4181.3,-17746.,-214.25,-21423.,-6491.2,-4586.8,-3126.2,82.637,2943.9,2684.4,2100.8,415.29,4599.1,1686.6,0.0000,7590.6,4449.7,4252.8,3658.0,0.0000,-517.03,-169.08,-114.38,-55.926,-193.26,-587.69,0.0000,-1100.2,-1654.3,-759.82,-1364.8
426.0000000000,113.67,2431.9,2538.6,2002.6,375.00,4193.2,974.40,0.98237,6369.4,2596.1,3350.1,1933.5,0.0000,-8957.5,-7752.0,-2061.3,-3006.2,-4176.9,-17742.,-213.88,-21420.,-6491.2,-4586.4,-3125.1,82.443,2937.0,2678.0,2091.1,414.23,4576.0,1686.6,0.0000,7576.6,4449.7,4252.8,3658.0,0.0000,-515.58,-168.54,-113.95,-55.786,-192.25,-587.69,0.0000,-1100.0,-1653.9,-759.82,-1364.3
427.0000000000,113.49,2427.5,2534.1,1998.9,374.21,4187.2,974.37,0.98328,6367.9,2596.4,3350.1,1934.0,0.0000,-8948.0,-7748.7,-2060.2,-3004.0,-4172.2,-17738.,-213.51,-21418.,-6491.1,-4586.1,-3124.0,82.317,2932.5,2673.9,2083.1,413.51,4556.8,1686.6,0.0000,7565.0,4449.7,4252.8,3658.0,0.0000,-514.55,-168.15,-113.61,-55.692,-191.40,-587.69,0.0000,-1099.8,-1653.6,-759.82,-1363.8
428.0000000000,113.38,2423.8,2530.4,1993.6,373.50,4178.9,974.37,0.98420,6365.4,2596.7,3350.1,1934.5,0.0000,-8938.5,-7745.4,-2059.0,-3001.8,-4167.2,-17734.,-213.13,-21415.,-6491.0,-4585.7,-3123.0,82.210,2928.7,2670.5,2075.7,412.90,4538.7,1686.6,0.0000,7554.0,4449.7,4252.8,3658.0,0.0000,-513.65,-167.79,-113.30,-55.612,-190.59,-587.69,0.0000,-1099.6,-1653.3,-759.81,-1363.4
429.0000000000,113.30,2420.4,2526.8,1987.2,372.82,4169.4,974.37,0.98511,6362.2,2597.1,3350.1,1935.0,0.0000,-8929.2,-7742.1,-2057.6,-2999.5,-4161.9,-17730.,-212.76,-21412.,-6490.9,-4585.4,-3121.9,82.032,2922.3,2664.7,2066.9,411.93,4517.8,1686.6,0.0000,7541.3,4449.7,4252.8,3658.0,0.0000,-512.30,-167.28,-112.91,-55.483,-189.67,-587.69,0.0000,-1099.4,-1653.0,-759.81,-1362.9
430.0000000000,113.13,2415.9,2522.1,1980.4,372.05,4158.6,974.37,0.98601,6357.8,2597.4,3350.1,1935.4,0.0000,-8919.7,-7738.7,-2056.1,-2997.3,-4156.5,-17726.,-212.39,-21409.,-6490.8,-4585.0,-3120.9,81.835,2915.3,2658.3,2057.7,410.86,4496.3,1686.6,0.0000,7528.3,4449.7,4252.8,3658.0,0.0000,-510.84,-166.74,-112.49,-55.342,-188.71,-587.69,0.0000,-1099.3,-1652.6,-759.81,-1362.4
431.0000000000,112.95,2411.1,2516.7,1973.0,371.18,4146.0,974.37,0.98691,6351.0,2597.7,3350.1,1935.9,0.0000,-8910.2,-7735.3,-2054.5,-2995.1,-4150.8,-17722.,-212.02,-21406.,-6490.6,-4584.6,-3119.9,81.638,2908.3,2651.9,2048.7,409.81,4474.9,1686.6,0.0000,7515.3,4449.7,4252.8,3658.0,0.0000,-509.38,-166.20,-112.08,-55.200,-187.76,-587.69,0.0000,-1099.1,-1652.3,-759.81,-1361.9
432.0000000000,112.75,2406.0,2511.4,1965.3,370.25,4130.7,974.36,0.98780,6342.4,2598.0,3350.1,1936.4,0.0000,-8900.6,-7731.8,-2052.7,-2992.8,-4144.9,-17718.,-211.65,-21403.,-6490.5,-4584.3,-3118.9,81.418,2900.5,2644.7,2039.1,408.63,4452.6,1686.6,0.0000,7501.8,4449.7,4252.8,3658.0,0.0000,-507.76,-165.61,-111.64,-55.043,-186.77,-587.69,0.0000,-1098.9,-1652.0,-759.81,-1361.5
433.0000000000,112.53,2400.5,2506.3,1957.1,369.31,4114.5,974.36,0.99961,6333.3,2598.4,3350.1,1936.8,0.0000,-8890.8,-7728.3,-2050.9,-2990.6,-4138.9,-17714.,-211.28,-21399.,-6490.4,-4583.9,-3117.9,81.242,2894.2,2639.0,2030.6,407.68,4432.5,1686.6,0.0000,7489.6,4449.7,4252.8,3658.0,0.0000,-506.43,-165.11,-111.26,-54.916,-185.87,-587.69,0.0000,-1098.7,-1651.7,-759.81,-1361.0
434.0000000000,112.33,2395.4,2500.9,1948.9,368.43,4098.5,974.36,1.0049,6323.7,2598.7,3350.1,1937.3,0.0000,-8881.1,-7724.8,-2049.0,-2988.3,-4132.6,-17711.,-210.92,-21396.,-6490.3,-4583.5,-3116.9,81.063,2887.8,2633.2,2022.1,406.71,4412.4,1686.6,0.0000,7477.4,4449.7,4252.8,3658.0,0.0000,-505.08,-164.61,-110.88,-54.786,-184.96,-587.69,0.0000,-1098.5,-1651.3,-759.81,-1360.5
435.0000000000,112.12,2390.3,2495.6,1940.9,367.55,4082.3,974.36,1.0058,6314.0,2599.0,3350.1,1937.8,0.0000,-8871.3,-7721.2,-2047.0,-2986.1,-4126.3,-17707.,-210.55,-21392.,-6490.2,-4583.1,-3115.9,80.854,2880.4,2626.4,2013.0,405.60,4391.1,1686.6,0.0000,7464.5,4449.7,4252.8,3658.0,0.0000,-503.54,-164.04,-110.46,-54.636,-184.01,-587.69,0.0000,-1098.3,-1651.0,-759.81,-1360.0
436.0000000000,111.91,2384.9,2489.8,1932.8,366.60,4065.4,974.36,1.0067,6303.9,2599.3,3350.1,1938.3,0.0000,-8861.4,-7717.6,-2045.0,-2983.8,-4119.8,-17703.,-210.19,-21389.,-6490.1,-4582.7,-3114.9,80.616,2871.9,2618.7,2003.3,404.34,4368.6,1686.6,0.0000,7450.9,4449.7,4252.8,3658.0,0.0000,-501.82,-163.42,-110.01,-54.467,-183.00,-587.69,0.0000,-1098.1,-1650.7,-759.81,-1359.6
437.0000000000,111.69,2379.1,2483.6,1924.6,365.62,4048.0,974.36,1.0076,6293.5,2599.6,3350.1,1938.7,0.0000,-8851.5,-7714.0,-2042.9,-2981.6,-4113.2,-17699.,-209.83,-21385.,-6489.9,-4582.3,-3114.0,80.437,2865.5,2612.9,1994.9,403.37,4348.7,1686.6,0.0000,7438.9,4449.7,4252.8,3658.0,0.0000,-500.47,-162.91,-109.62,-54.337,-182.11,-587.69,0.0000,-1097.9,-1650.4,-759.81,-1359.2
438.0000000000,111.48,2373.7,2477.7,1916.3,364.71,4030.4,974.35,1.0085,6283.2,2600.0,3350.1,1939.1,0.0000,-8841.5,-7710.4,-2040.8,-2979.3,-4106.4,-17695.,-209.47,-21381.,-6489.8,-4581.9,-3113.0,80.247,2858.8,2606.7,1986.3,402.35,4328.5,1686.6,0.0000,7426.6,4449.7,4252.8,3658.0,0.0000,-499.05,-162.38,-109.23,-54.200,-181.19,-587.69,0.0000,-1097.7,-1650.0,-759.81,-1358.7
439.0000000000,111.29,2368.2,2471.7,1908.0,363.77,4013.1,974.35,1.0094,6273.0,2600.3,3350.1,1939.6,0.0000,-8831.5,-7706.7,-2038.6,-2977.1,-4099.6,-17691.,-209.12,-21377.,-6489.7,-4581.5,-3112.0,80.014,2850.4,2599.1,1976.8,401.12,4306.5,1686.6,0.0000,7413.3,4449.7,4252.8,3658.0,0.0000,-497.36,-161.77,-108.79,-54.034,-180.20,-587.69,0.0000,-1097.5,-1649.7,-759.80,-1358.3
440.0000000000,110.88,2362.1,2465.3,1899.7,362.73,3995.7,974.32,1.0103,6262.5,2600.6,3350.1,1940.0,0.0000,-8821.4,-7703.0,-2036.3,-2974.8,-4092.6,-17687.,-208.77,-21373.,-6489.6,-4581.1,-3111.0,79.764,2841.6,2591.0,1967.0,399.81,4283.9,1686.6,0.0000,7399.5,4449.7,4252.8,3658.0,0.0000,-495.57,-161.12,-108.32,-53.857,-179.19,-587.69,0.0000,-1097.3,-1649.4,-759.80,-1357.9
441.0000000000,110.64,2355.9,2458.9,1891.2,361.70,3977.7,974.29,1.0175,6251.7,2600.9,3350.1,1940.5,0.0000,-8811.2,-7699.3,-2034.0,-2972.6,-4085.4,-17683.,-208.42,-21369.,-6489.4,-4580.7,-3110.1,79.587,2835.2,2585.3,1958.8,398.85,4264.5,1686.6,0.0000,7387.8,4449.7,4252.8,3658.0,0.0000,-494.23,-160.61,-107.95,-53.728,-178.31,-587.69,0.0000,-1097.2,-1649.1,-759.80,-1357.4
442.0000000000,110.43,2350.5,2453.0,1882.9,360.66,3959.9,974.27,1.0278,6241.0,2601.2,3350.1,1940.9,0.0000,-8801.0,-7695.6,-2031.7,-2970.3,-4078.1,-17679.,-208.08,-21365.,-6489.3,-4580.3,-3109.1,79.397,2828.5,2579.1,1950.3,397.84,4244.7,1686.6,0.0000,7375.8,4449.7,4252.8,3658.0,0.0000,-492.81,-160.09,-107.56,-53.591,-177.41,-587.69,0.0000,-1097.0,-1648.8,-759.80,-1357.0
443.0000000000,110.21,2344.9,2447.2,1874.7,359.71,3942.2,974.27,1.0287,6230.4,2601.6,3350.1,1941.3,0.0000,-8790.8,-7691.9,-2029.3,-2968.1,-4070.8,-17675.,-207.75,-21360.,-6489.2,-4579.9,-3108.1,79.153,2819.8,2571.2,1940.8,396.56,4222.8,1686.6,0.0000,7362.5,4449.7,4252.8,3658.0,0.0000,-491.06,-159.45,-107.11,-53.418,-176.42,-587.69,0.0000,-1096.8,-1648.4,-759.79,-1356.6
444.0000000000,109.99,2339.0,2441.0,1866.6,358.75,3924.5,974.26,1.0296,6219.3,2601.9,3350.1,1941.7,0.0000,-8780.5,-7688.1,-2026.9,-2965.8,-4063.3,-17671.,-207.42,-21356.,-6489.0,-4579.5,-3107.1,78.967,2813.1,2565.1,1932.5,395.56,4203.3,1686.6,0.0000,7350.7,4449.7,4252.8,3658.0,0.0000,-489.66,-158.93,-106.73,-53.284,-175.53,-587.69,0.0000,-1096.6,-1648.1,-759.79,-1356.2
445.0000000000,109.78,2333.3,2435.0,1858.5,357.80,3906.8,974.23,1.0345,6208.2,2602.2,3350.1,1942.2,0.0000,-8770.2,-7684.3,-2024.4,-2963.6,-4055.7,-17668.,-207.10,-21351.,-6488.9,-4579.1,-3106.2,78.755,2805.6,2558.2,1923.7,394.43,4182.9,1686.6,0.0000,7338.3,4449.7,4252.8,3658.0,0.0000,-488.11,-158.36,-106.32,-53.132,-174.61,-587.69,0.0000,-1096.4,-1647.8,-759.78,-1355.7
446.0000000000,109.55,2327.1,2428.6,1850.4,356.79,3888.8,974.21,1.0452,6196.9,2602.5,3350.1,1942.6,0.0000,-8759.9,-7680.6,-2021.9,-2961.3,-4048.1,-17664.,-206.78,-21347.,-6488.7,-4578.7,-3105.2,78.494,2796.3,2549.8,1914.0,393.07,4160.5,1686.6,0.0000,7324.8,4449.7,4252.8,3658.0,0.0000,-486.25,-157.69,-105.86,-52.947,-173.60,-587.69,0.0000,-1096.2,-1647.5,-759.78,-1355.3
447.0000000000,109.30,2320.6,2421.8,1842.0,355.72,3870.5,974.18,1.0461,6185.8,2602.8,3350.1,1943.0,0.0000,-8749.5,-7676.7,-2019.4,-2959.1,-4040.3,-17660.,-206.46,-21342.,-6488.6,-4578.2,-3104.2,78.267,2788.2,2542.4,1905.0,391.87,4139.6,1686.6,0.0000,7312.1,4449.7,4252.8,3658.0,0.0000,-484.60,-157.08,-105.43,-52.785,-172.65,-587.69,0.0000,-1096.0,-1647.2,-759.77,-1354.9
448.0000000000,109.07,2314.9,2415.8,1833.6,354.79,3852.4,974.18,1.0470,6174.7,2603.2,3350.1,1943.4,0.0000,-8739.1,-7672.9,-2016.8,-2956.8,-4032.4,-17656.,-206.14,-21337.,-6488.4,-4577.8,-3103.2,78.163,2784.5,2539.0,1898.2,391.28,4123.2,1686.6,0.0000,7302.2,4449.7,4252.8,3658.0,0.0000,-483.72,-156.73,-105.15,-52.707,-171.89,-587.69,0.0000,-1095.9,-1646.8,-759.77,-1354.5
449.0000000000,108.89,2310.1,2410.3,1825.7,353.95,3834.9,974.18,1.0479,6163.7,2603.5,3350.1,1943.8,0.0000,-8728.7,-7669.1,-2014.3,-2954.6,-4024.5,-17652.,-205.82,-21333.,-6488.3,-4577.4,-3102.2,77.944,2776.7,2531.9,1889.4,390.13,4102.9,1686.6,0.0000,7289.9,4449.7,4252.8,3658.0,0.0000,-482.13,-156.14,-104.73,-52.551,-170.96,-587.69,0.0000,-1095.7,-1646.5,-759.76,-1354.1
450.0000000000,108.67,2304.5,2404.3,1818.0,353.06,3817.3,974.18,1.0488,6152.8,2603.8,3350.1,1944.3,0.0000,-8718.3,-7665.3,-2011.7,-2952.4,-4016.5,-17648.,-205.50,-21328.,-6488.1,-4576.9,-3101.3,77.728,2769.0,2524.9,1880.7,388.98,4082.7,1686.6,0.0000,7277.6,4449.7,4252.8,3658.0,0.0000,-480.54,-155.56,-104.32,-52.396,-170.04,-587.69,0.0000,-1095.5,-1646.2,-759.76,-1353.6
451.0000000000,108.48,2298.7,2398.2,1810.0,352.14,3799.7,974.18,1.0496,6141.8,2604.2,3350.1,1944.7,0.0000,-8707.9,-7661.5,-2009.1,-2950.1,-4008.4,-17644.,-205.18,-21323.,-6487.9,-4576.5,-3100.3,77.522,2761.7,2518.2,1872.3,387.89,4063.2,1686.6,0.0000,7265.8,4449.7,4252.8,3658.0,0.0000,-479.03,-155.00,-103.93,-52.249,-169.16,-587.69,0.0000,-1095.3,-1645.9,-759.75,-1353.2
452.0000000000,108.25,2292.6,2391.7,1802.1,351.12,3781.7,974.18,1.0505,6130.7,2604.5,3350.1,1945.1,0.0000,-8697.5,-7657.7,-2006.4,-2947.9,-4000.3,-17640.,-204.87,-21318.,-6487.8,-4576.1,-3099.3,77.262,2752.4,2509.7,1862.8,386.54,4041.4,1686.6,0.0000,7252.6,4449.7,4252.8,3658.0,0.0000,-477.18,-154.34,-103.47,-52.065,-168.16,-587.69,0.0000,-1095.1,-1645.6,-759.75,-1352.8
453.0000000000,108.02,2285.9,2384.8,1794.0,350.04,3763.4,974.17,1.0514,6119.8,2604.8,3350.1,1945.5,0.0000,-8686.9,-7653.8,-2003.7,-2945.6,-3992.2,-17636.,-204.55,-21313.,-6487.6,-4575.6,-3098.3,77.016,2743.6,2501.7,1853.6,385.25,4020.3,1686.6,0.0000,7239.8,4449.7,4252.8,3658.0,0.0000,-475.42,-153.70,-103.03,-51.891,-167.20,-587.69,0.0000,-1094.9,-1645.3,-759.74,-1352.4
454.0000000000,107.91,2279.2,2377.9,1785.7,348.93,3745.2,974.17,1.0522,6108.9,2605.1,3350.1,1945.9,0.0000,-8676.3,-7649.9,-2001.0,-2943.4,-3983.9,-17632.,-204.24,-21308.,-6487.5,-4575.2,-3097.3,76.777,2735.1,2494.0,1844.6,384.00,3999.5,1686.6,0.0000,7227.2,4449.7,4252.8,3658.0,0.0000,-473.71,-153.07,-102.60,-51.721,-166.26,-587.69,0.0000,-1094.7,-1644.9,-759.74,-1352.0
455.0000000000,107.66,2272.6,2370.9,1777.2,347.81,3727.1,974.17,1.0531,6097.9,2605.4,3350.1,1946.3,0.0000,-8665.6,-7645.9,-1998.3,-2941.1,-3975.6,-17628.,-203.92,-21302.,-6487.3,-4574.7,-3096.3,76.526,2726.2,2485.9,1835.3,382.69,3978.2,1686.6,0.0000,7214.3,4449.7,4252.8,3658.0,0.0000,-471.92,-152.43,-102.15,-51.544,-165.29,-587.69,0.0000,-1094.6,-1644.6,-759.73,-1351.6
456.0000000000,107.40,2265.5,2363.7,1768.9,346.68,3708.7,974.17,1.0539,6086.7,2605.8,3350.1,1946.7,0.0000,-8654.8,-7642.0,-1995.5,-2938.8,-3967.3,-17624.,-203.61,-21297.,-6487.1,-4574.2,-3095.3,76.263,2716.8,2477.3,1825.8,381.32,3956.5,1686.6,0.0000,7201.2,4449.7,4252.8,3658.0,0.0000,-470.05,-151.75,-101.69,-51.357,-164.30,-587.69,0.0000,-1094.4,-1644.3,-759.73,-1351.2
457.0000000000,107.13,2258.1,2356.3,1760.4,345.51,3690.1,974.17,1.0548,6075.3,2606.1,3350.1,1947.1,0.0000,-8643.9,-7637.9,-1992.7,-2936.6,-3958.9,-17621.,-203.30,-21292.,-6486.9,-4573.8,-3094.3,75.994,2707.3,2468.6,1816.2,379.92,3934.7,1686.6,0.0000,7188.0,4449.7,4252.8,3658.0,0.0000,-468.15,-151.07,-101.22,-51.168,-163.31,-587.69,0.0000,-1094.2,-1644.0,-759.72,-1350.8
458.0000000000,106.86,2250.8,2348.7,1751.8,344.31,3671.2,974.17,1.0556,6063.7,2606.4,3350.1,1947.5,0.0000,-8633.0,-7633.9,-1989.8,-2934.3,-3950.5,-17617.,-202.99,-21286.,-6486.8,-4573.3,-3093.3,75.716,2697.3,2459.5,1806.5,378.48,3912.5,1686.6,0.0000,7174.6,4449.7,4252.8,3658.0,0.0000,-466.20,-150.36,-100.75,-50.972,-162.30,-587.69,0.0000,-1094.0,-1643.7,-759.72,-1350.4
459.0000000000,106.58,2244.3,2341.8,1743.3,343.27,3652.5,974.16,1.0565,6052.1,2606.7,3350.1,1947.9,0.0000,-8622.0,-7629.8,-1986.9,-2932.0,-3942.1,-17613.,-202.68,-21281.,-6486.6,-4572.8,-3092.4,75.631,2694.3,2456.8,1801.7,378.00,3900.9,1686.6,0.12086,7167.7,4449.8,4252.8,3658.0,0.0000,-465.43,-150.05,-100.54,-50.906,-161.74,-587.69,-0.55353E-02,-1093.8,-1643.4,-759.71,-1350.0
460.0000000000,106.40,2239.6,2336.1,1735.5,342.44,3635.2,974.16,1.0573,6040.8,2607.0,3350.1,1948.3,0.0000,-8611.1,-7625.8,-1984.1,-2929.8,-3933.8,-17609.,-202.37,-21275.,-6486.4,-4572.4,-3091.4,75.420,2686.8,2449.9,1793.4,376.89,3881.8,1686.6,0.0000,7156.0,4449.7,4252.8,3658.0,0.0000,-463.89,-149.48,-100.15,-50.755,-160.86,-587.69,0.0000,-1093.7,-1643.1,-759.70,-1349.6
461.0000000000,106.17,2234.1,2330.4,1728.1,341.47,3618.3,974.16,1.0581,6029.7,2607.3,3350.1,1948.8,0.0000,-8600.3,-7621.9,-1981.2,-2927.5,-3925.6,-17605.,-202.07,-21270.,-6486.2,-4571.9,-3090.4,75.214,2679.5,2443.2,1785.3,375.81,3863.1,1686.6,0.0000,7144.6,4449.7,4252.8,3658.0,0.0000,-462.38,-148.92,-99.764,-50.608,-160.00,-587.69,0.0000,-1093.5,-1642.8,-759.70,-1349.2
462.0000000000,105.99,2228.4,2324.2,1720.8,340.61,3601.1,974.16,1.0590,6018.5,2607.6,3350.1,1949.2,0.0000,-8589.4,-7617.9,-1978.4,-2925.3,-3917.5,-17601.,-201.76,-21264.,-6486.0,-4571.4,-3089.4,75.016,2672.4,2436.8,1777.3,374.76,3844.6,1686.6,0.0000,7133.4,4449.7,4252.8,3658.0,0.0000,-460.92,-148.38,-99.389,-50.466,-159.15,-587.69,0.0000,-1093.3,-1642.5,-759.69,-1348.8
463.0000000000,105.78,2222.7,2318.1,1713.3,339.72,3584.0,974.16,1.0598,6007.4,2607.8,3350.1,1949.6,0.0000,-8578.6,-7613.9,-1975.5,-2923.1,-3909.5,-17597.,-201.46,-21259.,-6485.9,-4570.9,-3088.4,74.845,2666.3,2431.2,1769.9,373.85,3827.3,1686.6,0.0000,7122.9,4449.7,4252.8,3658.0,0.0000,-459.63,-147.92,-99.048,-50.343,-158.34,-587.69,0.0000,-1093.1,-1642.2,-759.69,-1348.4
464.0000000000,105.58,2217.3,2312.2,1706.0,338.85,3566.8,974.16,1.0606,5996.7,2608.1,3350.1,1950.0,0.0000,-8567.9,-7609.9,-1972.6,-2920.8,-3901.6,-17593.,-201.16,-21253.,-6485.7,-4570.5,-3087.4,74.638,2658.9,2424.5,1761.8,372.76,3808.6,1686.6,0.0000,7111.6,4449.7,4252.8,3658.0,0.0000,-458.12,-147.39,-98.665,-50.196,-157.48,-587.69,0.0000,-1093.0,-1641.9,-759.68,-1348.0
465.0000000000,105.37,2211.4,2306.2,1698.4,337.93,3550.1,974.15,1.0615,5986.6,2608.4,3350.1,1950.3,0.0000,-8557.1,-7605.9,-1969.7,-2918.6,-3893.9,-17589.,-200.87,-21247.,-6485.5,-4570.0,-3086.4,74.407,2650.7,2417.0,1753.3,371.56,3789.0,1686.6,0.0000,7099.7,4449.7,4252.8,3658.0,0.0000,-456.46,-146.82,-98.254,-50.032,-156.57,-587.69,0.0000,-1092.8,-1641.6,-759.67,-1347.6
466.0000000000,105.28,2205.1,2300.2,1690.7,336.92,3533.6,974.15,1.0623,5976.5,2608.7,3350.0,1950.7,0.0000,-8546.2,-7602.0,-1966.8,-2916.4,-3886.3,-17585.,-200.58,-21241.,-6485.3,-4569.5,-3085.4,74.151,2641.6,2408.7,1744.3,370.23,3768.5,1686.6,0.0000,7087.3,4449.7,4252.8,3658.0,0.0000,-454.65,-146.19,-97.814,-49.851,-155.63,-587.69,0.0000,-1092.6,-1641.4,-759.67,-1347.2
467.0000000000,105.09,2198.4,2293.3,1682.9,335.82,3516.6,974.09,1.0631,5966.1,2609.0,3350.0,1951.1,0.0000,-8535.4,-7598.0,-1963.9,-2914.1,-3879.0,-17581.,-200.29,-21236.,-6485.1,-4569.0,-3084.4,73.899,2632.6,2400.5,1735.4,368.92,3748.3,1686.6,0.0000,7075.1,4449.7,4252.8,3658.0,0.0000,-452.86,-145.58,-97.380,-49.674,-154.70,-587.69,0.0000,-1092.4,-1641.1,-759.66,-1346.9
468.0000000000,104.83,2191.5,2286.1,1674.9,334.70,3499.2,974.08,1.0639,5955.6,2609.3,3350.0,1951.5,0.0000,-8524.4,-7593.9,-1960.9,-2911.9,-3871.7,-17577.,-199.99,-21230.,-6484.9,-4568.5,-3083.4,73.644,2623.5,2392.2,1726.5,367.60,3728.0,1686.6,0.0000,7062.8,4449.7,4252.8,3658.0,0.0000,-451.06,-144.96,-96.944,-49.494,-153.76,-587.69,0.0000,-1092.2,-1640.8,-759.65,-1346.5
469.0000000000,104.57,2184.8,2279.0,1666.8,333.60,3481.7,974.08,1.0647,5945.0,2609.6,3350.0,1951.9,0.0000,-8513.4,-7589.8,-1957.9,-2909.6,-3864.6,-17573.,-199.70,-21224.,-6484.7,-4568.0,-3082.4,73.428,2615.8,2385.2,1718.2,366.46,3709.1,1686.6,0.0000,7051.3,4449.7,4252.8,3658.0,0.0000,-449.50,-144.41,-96.551,-49.340,-152.87,-587.69,0.0000,-1092.1,-1640.5,-759.64,-1346.1
470.0000000000,104.33,2178.7,2272.4,1658.8,332.63,3464.5,974.07,1.0655,5934.4,2609.9,3350.1,1952.3,0.0000,-8502.4,-7585.8,-1954.9,-2907.4,-3857.4,-17569.,-199.41,-21218.,-6484.5,-4567.5,-3081.4,73.278,2610.5,2380.3,1711.5,365.66,3693.2,1686.6,0.0000,7041.7,4449.7,4252.8,3658.0,0.0000,-448.34,-144.00,-96.242,-49.231,-152.09,-587.69,0.0000,-1091.9,-1640.2,-759.64,-1345.7
471.0000000000,104.12,2173.5,2266.7,1651.1,331.80,3448.0,974.05,1.0663,5923.9,2610.1,3350.1,1952.7,0.0000,-8491.5,-7581.8,-1951.9,-2905.2,-3850.3,-17565.,-199.13,-21212.,-6484.3,-4566.9,-3080.4,73.117,2604.7,2375.1,1704.5,364.80,3676.9,1686.6,0.0000,7031.8,4449.7,4252.8,3658.0,0.0000,-447.12,-143.56,-95.921,-49.115,-151.29,-587.69,0.0000,-1091.7,-1639.9,-759.63,-1345.3
472.0000000000,103.78,2168.4,2261.3,1644.0,331.00,3431.8,974.05,1.0671,5913.3,2610.4,3350.1,1953.0,0.0000,-8480.6,-7577.9,-1948.9,-2903.0,-3843.1,-17561.,-198.84,-21206.,-6484.1,-4566.4,-3079.4,72.916,2597.6,2368.6,1696.8,363.75,3659.1,1686.6,0.0000,7021.1,4449.7,4252.8,3658.0,0.0000,-445.65,-143.05,-95.554,-48.972,-150.43,-587.69,0.0000,-1091.6,-1639.6,-759.62,-1345.0
473.0000000000,103.58,2162.7,2255.4,1636.8,330.16,3415.5,974.04,1.0679,5902.6,2610.7,3350.1,1953.4,0.0000,-8469.8,-7574.0,-1945.9,-2900.8,-3835.9,-17558.,-198.55,-21200.,-6483.9,-4565.9,-3078.4,72.691,2589.6,2361.3,1688.6,362.58,3640.4,1686.6,0.0000,7009.7,4449.7,4252.8,3658.0,0.0000,-444.04,-142.50,-95.159,-48.813,-149.52,-587.69,0.0000,-1091.4,-1639.4,-759.61,-1344.6
474.0000000000,103.37,2156.6,2249.0,1629.4,329.21,3398.9,974.04,1.0687,5892.0,2611.0,3350.1,1953.8,0.0000,-8458.9,-7570.0,-1942.9,-2898.5,-3828.7,-17554.,-198.26,-21194.,-6483.7,-4565.4,-3077.4,72.460,2581.3,2353.7,1680.4,361.37,3621.5,1686.6,0.0000,6998.3,4449.7,4252.8,3658.0,0.0000,-442.39,-141.93,-94.756,-48.649,-148.61,-587.69,0.0000,-1091.2,-1639.1,-759.61,-1344.2
475.0000000000,103.14,2150.5,2242.5,1621.9,328.22,3382.2,974.02,1.0695,5881.8,2611.3,3350.1,1954.2,0.0000,-8448.0,-7566.1,-1939.9,-2896.3,-3821.5,-17550.,-197.98,-21187.,-6483.5,-4564.9,-3076.5,72.260,2574.2,2347.3,1672.7,360.32,3604.0,1686.6,0.0000,6987.6,4449.7,4252.8,3658.0,0.0000,-440.93,-141.42,-94.392,-48.507,-147.75,-587.69,0.0000,-1091.0,-1638.8,-759.60,-1343.8
476.0000000000,102.92,2144.4,2236.2,1614.4,327.25,3365.8,973.99,1.0703,5871.7,2611.6,3350.1,1954.5,0.0000,-8437.2,-7562.1,-1936.9,-2894.1,-3814.2,-17546.,-197.69,-21181.,-6483.2,-4564.3,-3075.5,72.037,2566.3,2340.0,1664.7,359.16,3585.6,1686.6,0.0000,6976.5,4449.7,4252.8,3658.0,0.0000,-439.34,-140.87,-94.003,-48.350,-146.86,-587.69,0.0000,-1090.9,-1638.5,-759.59,-1343.5
477.0000000000,102.68,2138.2,2229.7,1606.9,326.24,3349.7,974.01,1.0711,5861.8,2611.8,3350.1,1954.9,0.0000,-8426.3,-7558.1,-1933.8,-2891.9,-3806.9,-17542.,-197.41,-21175.,-6483.0,-4563.8,-3074.5,71.789,2557.5,2332.0,1656.2,357.88,3566.3,1686.6,0.0000,6964.8,4449.7,4252.8,3658.0,0.0000,-437.59,-140.27,-93.584,-48.175,-145.93,-587.69,0.0000,-1090.7,-1638.2,-759.58,-1343.1
478.0000000000,102.44,2131.6,2222.7,1599.2,325.17,3333.5,974.03,1.0719,5851.7,2612.1,3350.1,1955.3,0.0000,-8415.3,-7554.1,-1930.8,-2889.7,-3799.6,-17538.,-197.12,-21169.,-6482.8,-4563.3,-3073.5,71.538,2548.5,2323.8,1647.6,356.58,3546.9,1686.6,0.0000,6953.1,4449.7,4252.8,3658.0,0.0000,-435.82,-139.66,-93.161,-47.998,-144.99,-587.69,0.0000,-1090.5,-1637.9,-759.58,-1342.7
479.0000000000,102.19,2124.7,2215.5,1591.5,324.06,3316.9,974.03,1.0727,5841.6,2612.4,3350.1,1955.7,0.0000,-8404.4,-7550.1,-1927.7,-2887.5,-3792.2,-17534.,-196.84,-21163.,-6482.6,-4562.7,-3072.5,71.280,2539.3,2315.4,1639.0,355.25,3527.3,1686.6,0.0000,6941.2,4449.7,4252.8,3658.0,0.0000,-434.02,-139.04,-92.733,-47.817,-144.04,-587.69,0.0000,-1090.3,-1637.7,-759.57,-1342.3
480.0000000000,101.93,2117.9,2208.2,1583.7,322.92,3300.1,974.02,1.0734,5831.3,2612.7,3350.1,1956.0,0.0000,-8393.3,-7546.0,-1924.5,-2885.2,-3784.8,-17530.,-196.56,-21156.,-6482.4,-4562.2,-3071.5,71.044,2530.9,2307.8,1630.7,354.02,3508.6,1686.6,0.0000,6929.9,4449.7,4252.8,3658.0,0.0000,-432.34,-138.46,-92.330,-47.651,-143.13,-587.69,0.0000,-1090.1,-1637.4,-759.56,-1342.0
481.0000000000,101.68,2111.3,2201.1,1575.8,321.83,3283.2,974.00,1.0742,5820.9,2613.0,3350.1,1956.4,0.0000,-8382.3,-7542.0,-1921.4,-2883.0,-3777.3,-17526.,-196.27,-21150.,-6482.1,-4561.6,-3070.5,70.800,2522.2,2299.9,1622.4,352.76,3489.7,1686.6,0.0000,6918.4,4449.7,4252.8,3658.0,0.0000,-430.62,-137.87,-91.919,-47.479,-142.21,-587.69,0.0000,-1090.0,-1637.1,-759.55,-1341.6
482.0000000000,101.43,2104.5,2193.8,1567.9,320.72,3266.4,974.00,1.0750,5810.7,2613.2,3350.1,1956.8,0.0000,-8371.2,-7537.9,-1918.2,-2880.8,-3769.9,-17522.,-195.99,-21143.,-6481.9,-4561.1,-3069.5,70.543,2513.0,2291.5,1613.8,351.43,3470.3,1686.6,0.0000,6906.7,4449.7,4252.8,3658.0,0.0000,-428.82,-137.25,-91.493,-47.298,-141.27,-587.69,0.0000,-1089.8,-1636.8,-759.54,-1341.3
483.0000000000,101.18,2097.5,2186.5,1560.0,319.61,3249.5,974.00,1.0757,5800.3,2613.5,3350.2,1957.1,0.0000,-8360.1,-7533.8,-1915.1,-2878.6,-3762.4,-17518.,-195.72,-21137.,-6481.7,-4560.5,-3068.5,70.295,2504.2,2283.4,1605.4,350.15,3451.3,1686.6,0.0000,6895.2,4449.7,4252.8,3658.0,0.0000,-427.08,-136.65,-91.079,-47.124,-140.35,-587.69,0.0000,-1089.6,-1636.6,-759.53,-1340.9
484.0000000000,100.92,2090.6,2179.3,1552.2,318.52,3232.6,974.00,1.0765,5789.7,2613.7,3350.2,1957.5,0.0000,-8349.0,-7529.7,-1911.9,-2876.3,-3754.8,-17514.,-195.44,-21130.,-6481.4,-4560.0,-3067.5,70.060,2495.9,2275.8,1597.4,348.93,3433.0,1686.6,0.0000,6884.1,4449.7,4252.8,3658.0,0.0000,-425.41,-136.08,-90.681,-46.958,-139.45,-587.69,0.0000,-1089.4,-1636.4,-759.52,-1340.5
485.0000000000,100.67,2084.1,2172.4,1544.4,317.47,3215.8,974.00,1.0773,5779.2,2614.0,3350.2,1957.9,0.0000,-8337.9,-7525.5,-1908.7,-2874.1,-3747.3,-17510.,-195.17,-21124.,-6481.2,-4559.4,-3066.5,69.860,2488.7,2269.3,1590.0,347.89,3416.1,1686.6,0.0000,6873.9,4449.7,4252.8,3658.0,0.0000,-423.96,-135.57,-90.326,-46.816,-138.62,-587.69,0.0000,-1089.3,-1636.1,-759.52,-1340.2
486.0000000000,100.44,2078.2,2166.1,1536.8,316.54,3199.3,973.98,1.0780,5768.7,2614.2,3350.2,1958.2,0.0000,-8326.9,-7521.4,-1905.5,-2871.9,-3739.7,-17506.,-194.89,-21117.,-6481.0,-4558.9,-3065.5,69.690,2482.7,2263.8,1583.2,346.99,3400.4,1686.6,0.0000,6864.4,4449.7,4252.8,3658.0,0.0000,-422.69,-135.13,-90.007,-46.694,-137.83,-587.69,0.0000,-1089.1,-1635.9,-759.51,-1339.8
487.0000000000,100.24,2072.8,2160.5,1529.5,315.70,3183.4,973.96,1.0788,5758.5,2614.4,3350.2,1958.5,0.0000,-8316.0,-7517.4,-1902.3,-2869.7,-3732.1,-17502.,-194.63,-21111.,-6480.7,-4558.3,-3064.5,69.524,2476.8,2258.4,1576.6,346.12,3385.0,1686.6,0.0000,6855.1,4449.7,4252.8,3658.0,0.0000,-421.45,-134.69,-89.694,-46.575,-137.05,-587.69,0.0000,-1089.0,-1635.7,-759.50,-1339.5
488.0000000000,100.04,2067.7,2154.5,1522.6,314.93,3167.9,973.96,1.0795,5748.3,2614.7,3350.2,1958.9,0.0000,-8305.2,-7513.4,-1899.1,-2867.5,-3724.6,-17498.,-194.36,-21104.,-6480.5,-4557.7,-3063.5,69.351,2470.6,2252.8,1569.8,345.21,3369.4,1686.6,0.0000,6845.6,4449.7,4252.8,3658.0,0.0000,-420.16,-134.24,-89.374,-46.452,-136.27,-587.69,0.0000,-1088.8,-1635.4,-759.49,-1339.2
489.0000000000,99.859,2062.5,2148.9,1515.8,314.13,3152.6,973.95,1.0803,5738.3,2614.9,3350.2,1959.2,0.0000,-8294.4,-7509.4,-1895.9,-2865.3,-3717.0,-17494.,-194.10,-21098.,-6480.3,-4557.2,-3062.5,69.158,2463.7,2246.5,1562.7,344.20,3353.1,1686.6,0.0000,6835.7,4449.7,4252.8,3658.0,0.0000,-418.76,-133.76,-89.031,-46.315,-135.45,-587.69,0.0000,-1088.6,-1635.2,-759.48,-1338.9
490.0000000000,99.665,2056.9,2143.0,1509.1,313.27,3137.3,973.95,1.0810,5728.5,2615.1,3350.2,1959.5,0.0000,-8283.7,-7505.5,-1892.7,-2863.1,-3709.5,-17490.,-193.84,-21091.,-6480.0,-4556.6,-3061.5,68.936,2455.8,2239.3,1555.0,343.05,3335.6,1686.6,0.0000,6825.2,4449.7,4252.8,3658.0,0.0000,-417.18,-133.22,-88.654,-46.159,-134.59,-587.69,0.0000,-1088.5,-1634.9,-759.47,-1338.5
491.0000000000,99.452,2050.9,2137.0,1502.2,312.33,3121.9,973.95,1.0818,5718.8,2615.4,3350.2,1959.9,0.0000,-8272.9,-7501.5,-1889.6,-2860.9,-3701.9,-17486.,-193.58,-21085.,-6479.8,-4556.0,-3060.5,68.703,2447.5,2231.7,1547.1,341.84,3317.8,1686.6,0.0000,6814.4,4449.7,4252.8,3658.0,0.0000,-415.52,-132.65,-88.265,-45.995,-133.72,-587.69,0.0000,-1088.3,-1634.7,-759.46,-1338.2
492.0000000000,99.199,2045.8,2131.6,1495.3,311.54,3106.5,973.95,1.0825,5709.4,2615.6,3350.2,1960.2,0.0000,-8262.2,-7497.6,-1886.4,-2858.7,-3694.3,-17483.,-193.33,-21078.,-6479.5,-4555.4,-3059.5,68.718,2448.1,2232.2,1543.8,341.86,3308.8,1686.6,0.0000,6808.8,4449.7,4252.8,3658.0,0.0000,-415.37,-132.57,-88.155,-45.998,-133.20,-587.69,0.0000,-1088.2,-1634.5,-759.45,-1337.9
493.0000000000,98.972,2042.4,2127.6,1488.8,310.96,3092.3,973.92,1.0833,5700.3,2615.9,3350.2,1960.5,0.0000,-8251.7,-7493.7,-1883.3,-2856.6,-3686.7,-17479.,-193.07,-21071.,-6479.3,-4554.9,-3058.5,68.490,2439.9,2224.8,1536.0,340.68,3291.3,1686.6,0.0000,6798.3,4449.7,4252.8,3658.0,0.0000,-413.75,-132.02,-87.774,-45.838,-132.34,-587.69,0.0000,-1088.0,-1634.2,-759.44,-1337.5
494.0000000000,98.762,2037.7,2122.9,1482.7,310.16,3078.2,973.90,1.0840,5691.5,2616.1,3350.2,1960.9,0.0000,-8241.2,-7489.9,-1880.1,-2854.4,-3679.1,-17475.,-192.82,-21065.,-6479.0,-4554.3,-3057.5,68.340,2434.6,2219.9,1528.8,339.86,3274.3,1686.6,0.0000,6788.0,4449.7,4252.8,3658.0,0.0000,-412.61,-131.62,-87.451,-45.730,-131.50,-587.69,0.0000,-1087.8,-1634.0,-759.43,-1337.2
495.0000000000,98.628,2034.0,2118.5,1476.3,309.70,3064.0,973.85,0.92112,5682.6,2616.3,3350.2,1961.2,0.0000,-8230.9,-7486.2,-1877.0,-2852.2,-3671.5,-17471.,-192.56,-21058.,-6478.8,-4553.7,-3056.5,68.386,2435.6,2220.9,1524.5,339.92,3262.7,1686.6,0.0000,6780.9,4449.7,4252.8,3658.0,0.0000,-412.54,-131.57,-87.316,-45.742,-130.88,-587.69,0.0000,-1087.7,-1633.8,-759.42,-1336.9
496.0000000000,98.558,2031.3,2115.3,1470.2,309.19,3050.1,973.83,0.89248,5673.5,2616.6,3350.2,1961.5,0.0000,-8220.7,-7482.5,-1873.8,-2850.1,-3663.8,-17467.,-192.31,-21051.,-6478.5,-4553.1,-3055.5,68.149,2427.8,2213.7,1517.0,338.78,3245.7,1686.6,0.0000,6770.6,4449.7,4252.8,3658.0,0.0000,-410.98,-131.04,-86.947,-45.589,-130.03,-587.69,0.0000,-1087.5,-1633.5,-759.41,-1336.6
497.0000000000,98.371,2026.8,2110.7,1464.2,308.44,3035.9,973.83,0.89309,5664.6,2616.8,3350.2,1961.8,0.0000,-8210.5,-7478.9,-1870.7,-2848.0,-3656.2,-17463.,-192.05,-21045.,-6478.3,-4552.5,-3054.5,67.940,2420.3,2206.9,1509.6,337.70,3228.8,1686.6,0.0000,6760.4,4449.7,4252.8,3658.0,0.0000,-409.49,-130.53,-86.586,-45.442,-129.20,-587.69,0.0000,-1087.4,-1633.3,-759.40,-1336.2
498.0000000000,98.221,2023.2,2106.7,1458.0,308.01,3021.6,973.83,0.89370,5655.8,2617.0,3350.3,1962.2,0.0000,-8200.4,-7475.3,-1867.6,-2845.9,-3648.6,-17459.,-191.80,-21038.,-6478.0,-4551.9,-3053.5,68.156,2425.7,2211.9,1507.5,338.34,3221.7,1686.6,0.0000,6756.1,4449.7,4252.8,3658.0,0.0000,-410.12,-130.71,-86.587,-45.531,-128.76,-587.69,0.0000,-1087.3,-1633.1,-759.39,-1335.9
499.0000000000,98.216,2022.7,2105.8,1452.1,307.86,3008.7,973.83,0.89430,5647.5,2617.3,3350.3,1962.5,0.0000,-8190.6,-7471.9,-1864.5,-2843.8,-3641.0,-17455.,-191.54,-21031.,-6477.8,-4551.3,-3052.5,68.068,2424.9,2211.1,1503.1,338.18,3210.7,1686.6,0.0000,6749.4,4449.7,4252.8,3658.0,0.0000,-409.80,-130.58,-86.432,-45.515,-128.17,-587.69,0.0000,-1087.1,-1632.9,-759.38,-1335.6
500.0000000000,98.140,2021.7,2104.4,1447.1,307.58,2996.7,973.83,0.89490,5639.4,2617.5,3350.3,1962.8,0.0000,-8181.1,-7468.6,-1861.4,-2841.7,-3633.4,-17451.,-191.29,-21024.,-6477.5,-4550.7,-3051.5,67.945,2420.5,2207.1,1497.4,337.51,3197.0,1686.6,0.0000,6741.1,4449.7,4252.8,3658.0,0.0000,-408.83,-130.24,-86.170,-45.426,-127.46,-587.69,0.0000,-1087.0,-1632.6,-759.37,-1335.3
501.0000000000,98.067,2019.0,2101.4,1442.2,307.28,2984.3,973.83,0.89549,5631.2,2617.7,3350.3,1963.1,0.0000,-8171.6,-7465.3,-1858.4,-2839.7,-3625.9,-17447.,-191.04,-21018.,-6477.2,-4550.1,-3050.5,67.792,2415.0,2202.1,1491.1,336.70,3182.5,1686.6,0.0000,6732.3,4449.7,4252.8,3658.0,0.0000,-407.69,-129.85,-85.878,-45.318,-126.73,-587.69,0.0000,-1086.9,-1632.4,-759.36,-1335.0
502.0000000000,97.969,2015.1,2097.6,1437.0,306.68,2971.6,973.80,0.89608,5623.1,2617.9,3350.3,1963.5,0.0000,-8162.2,-7462.0,-1855.3,-2837.6,-3618.3,-17443.,-190.78,-21011.,-6477.0,-4549.5,-3049.5,67.595,2408.0,2195.7,1484.1,335.68,3166.7,1686.6,0.0000,6722.7,4449.7,4252.8,3658.0,0.0000,-406.28,-129.38,-85.538,-45.180,-125.94,-587.69,0.0000,-1086.7,-1632.2,-759.35,-1334.7
503.0000000000,97.803,2010.7,2092.8,1431.3,305.88,2958.4,973.78,0.89667,5614.9,2618.2,3350.3,1963.8,0.0000,-8152.6,-7458.7,-1852.2,-2835.6,-3610.7,-17439.,-190.53,-21004.,-6476.7,-4548.9,-3048.5,67.392,2400.8,2189.1,1477.1,334.63,3150.7,1686.6,0.0000,6713.0,4449.7,4252.8,3658.0,0.0000,-404.84,-128.89,-85.194,-45.037,-125.14,-587.69,0.0000,-1086.5,-1631.9,-759.34,-1334.3
504.0000000000,97.610,2005.5,2087.4,1425.5,305.04,2944.7,973.78,0.89725,5606.5,2618.4,3350.4,1964.1,0.0000,-8143.0,-7455.3,-1849.2,-2833.5,-3603.1,-17435.,-190.28,-20998.,-6476.5,-4548.3,-3047.5,67.195,2393.8,2182.7,1470.3,333.61,3135.2,1686.6,0.0000,6703.6,4449.7,4252.8,3658.0,0.0000,-403.44,-128.42,-84.858,-44.899,-124.37,-587.69,0.0000,-1086.4,-1631.7,-759.33,-1334.0
505.0000000000,97.407,2000.3,2082.0,1419.3,304.15,2931.3,973.78,0.89785,5598.7,2618.6,3350.4,1964.4,0.0000,-8133.3,-7451.9,-1846.1,-2831.4,-3595.5,-17431.,-190.03,-20991.,-6476.2,-4547.6,-3046.5,66.991,2386.5,2176.1,1463.3,332.55,3119.4,1686.6,0.0000,6694.1,4449.7,4252.8,3658.0,0.0000,-401.99,-127.93,-84.516,-44.756,-123.58,-587.69,0.0000,-1086.2,-1631.5,-759.32,-1333.7
506.0000000000,97.299,1995.4,2076.7,1412.8,303.25,2918.2,973.76,0.89843,5591.2,2618.9,3350.4,1964.7,0.0000,-8123.6,-7448.4,-1842.9,-2829.3,-3587.8,-17427.,-189.78,-20984.,-6475.9,-4547.0,-3045.5,66.788,2379.3,2169.5,1456.5,331.50,3103.9,1686.6,0.0000,6684.7,4449.7,4252.8,3658.0,0.0000,-400.55,-127.44,-84.177,-44.614,-122.81,-587.69,0.0000,-1086.1,-1631.2,-759.31,-1333.4
507.0000000000,97.174,1989.8,2071.1,1406.6,302.34,2905.2,973.76,0.89901,5583.2,2619.1,3350.4,1965.1,0.0000,-8113.8,-7444.9,-1839.8,-2827.2,-3580.1,-17423.,-189.53,-20977.,-6475.6,-4546.4,-3044.4,66.574,2371.7,2162.6,1449.5,330.40,3088.0,1686.6,0.0000,6675.1,4449.7,4252.8,3658.0,0.0000,-399.05,-126.94,-83.826,-44.464,-122.02,-587.69,0.0000,-1085.9,-1631.0,-759.30,-1333.1
508.0000000000,96.957,1984.5,2065.5,1400.3,301.45,2891.9,973.76,0.89959,5575.0,2619.3,3350.5,1965.4,0.0000,-8103.9,-7441.4,-1836.7,-2825.1,-3572.4,-17419.,-189.28,-20970.,-6475.4,-4545.8,-3043.4,66.419,2366.2,2157.5,1443.8,329.59,3075.1,1686.6,0.0000,6667.3,4449.7,4252.8,3658.0,0.0000,-397.90,-126.54,-83.554,-44.354,-121.35,-587.69,0.0000,-1085.8,-1630.8,-759.28,-1332.8
509.0000000000,96.768,1979.6,2060.2,1394.1,300.63,2878.5,973.75,0.90017,5566.7,2619.5,3350.5,1965.7,0.0000,-8094.1,-7437.9,-1833.5,-2823.1,-3564.7,-17415.,-189.03,-20964.,-6475.1,-4545.1,-3042.4,66.217,2358.9,2151.0,1437.0,328.55,3059.8,1686.6,0.0000,6658.0,4449.7,4252.8,3658.0,0.0000,-396.47,-126.06,-83.218,-44.212,-120.58,-587.69,0.0000,-1085.6,-1630.6,-759.27,-1332.5
510.0000000000,96.447,1974.9,2055.2,1388.2,299.85,2865.2,973.73,0.90071,5558.3,2619.8,3350.5,1966.0,0.0000,-8084.2,-7434.5,-1830.3,-2821.0,-3557.0,-17412.,-188.78,-20957.,-6474.8,-4544.5,-3041.4,66.132,2355.9,2148.2,1434.0,328.11,3052.9,1686.6,0.0000,6653.8,4449.7,4252.8,3658.0,0.0000,-395.74,-125.80,-83.069,-44.149,-120.16,-587.69,0.0000,-1085.5,-1630.3,-759.26,-1332.2
511.0000000000,96.307,1978.8,2057.9,1383.1,300.65,2854.2,973.72,0.90130,5550.3,2620.0,3350.5,1966.3,0.0000,-8075.1,-7431.4,-1827.4,-2819.0,-3549.4,-17408.,-188.53,-20950.,-6474.5,-4543.9,-3040.4,69.379,2411.2,2198.4,1453.6,335.55,3087.1,1686.6,0.63312,6674.2,4450.0,4253.1,3658.3,0.0000,-404.33,-128.56,-84.484,-45.128,-121.36,-587.69,-0.28998E-01,-1085.7,-1630.1,-759.25,-1331.9
512.0000000000,97.015,1997.1,2072.5,1381.4,303.51,2848.3,973.70,0.90189,5543.8,2620.2,3350.5,1943.3,0.0000,-8067.8,-7429.2,-1824.6,-2817.2,-3542.0,-17404.,-188.29,-20943.,-6474.3,-4543.2,-3039.5,68.139,2427.4,2213.4,1453.0,337.65,3079.4,1686.6,0.0000,6669.5,4449.7,4252.8,3658.0,0.0000,-407.36,-129.46,-84.748,-45.482,-120.92,-587.69,0.0000,-1085.6,-1629.9,-759.24,-1331.6
513.0000000000,97.420,2010.5,2086.1,1382.7,305.29,2843.7,973.70,0.90246,5538.1,2620.4,3350.5,1943.6,0.0000,-8061.4,-7427.7,-1821.9,-2815.5,-3534.9,-17400.,-188.05,-20937.,-6474.0,-4542.6,-3038.5,68.169,2428.5,2214.4,1447.6,337.69,3065.1,1686.6,0.0000,6660.8,4449.7,4252.8,3658.0,0.0000,-407.35,-129.45,-84.580,-45.499,-120.20,-587.69,0.0000,-1085.4,-1629.7,-759.23,-1331.2
514.0000000000,97.777,2015.7,2091.4,1382.4,306.84,2836.7,973.70,0.90306,5532.3,2620.7,3350.5,1943.9,0.0000,-8055.2,-7426.1,-1819.3,-2813.8,-3527.8,-17396.,-187.80,-20930.,-6473.7,-4542.0,-3037.4,68.098,2426.0,2212.1,1441.7,337.26,3050.7,1686.6,0.0000,6652.0,4449.7,4252.8,3658.0,0.0000,-406.75,-129.25,-84.343,-45.449,-119.48,-587.69,0.0000,-1085.3,-1629.5,-759.22,-1330.9
515.0000000000,98.035,2016.2,2093.3,1380.8,307.00,2827.6,973.67,0.90362,5525.9,2620.9,3350.6,1944.2,0.0000,-8049.0,-7424.4,-1816.6,-2812.0,-3520.7,-17392.,-187.56,-20924.,-6473.4,-4541.3,-3036.4,67.969,2421.4,2207.9,1435.5,336.56,3035.9,1686.6,0.0000,6643.1,4449.7,4252.8,3658.0,0.0000,-405.81,-128.93,-84.063,-45.359,-118.74,-587.69,0.0000,-1085.1,-1629.2,-759.20,-1330.6
516.0000000000,98.013,2014.7,2092.1,1377.3,306.52,2817.3,973.62,0.90417,5520.0,2621.1,3350.6,1944.5,0.0000,-8042.5,-7422.6,-1814.0,-2810.2,-3513.4,-17388.,-187.31,-20917.,-6473.1,-4540.7,-3035.4,67.800,2415.3,2202.4,1428.9,335.67,3020.8,1686.6,0.0000,6633.9,4449.7,4252.8,3658.0,0.0000,-404.63,-128.54,-83.751,-45.242,-118.00,-587.69,0.0000,-1085.0,-1629.0,-759.19,-1330.3
517.0000000000,97.881,2012.0,2089.7,1373.2,305.86,2806.0,973.62,0.91375,5514.5,2621.3,3350.6,1944.7,0.0000,-8035.7,-7420.5,-1811.3,-2808.4,-3506.1,-17384.,-187.06,-20910.,-6472.9,-4540.0,-3034.4,67.638,2409.6,2197.1,1422.8,334.83,3006.7,1686.6,0.0000,6625.4,4449.7,4252.8,3658.0,0.0000,-403.50,-128.17,-83.458,-45.129,-117.29,-587.69,0.0000,-1084.8,-1628.8,-759.18,-1330.1
518.0000000000,97.726,2008.4,2087.2,1367.8,305.11,2796.3,973.62,0.91846,5511.7,2621.6,3350.6,1945.0,0.0000,-8028.8,-7418.4,-1808.5,-2806.5,-3498.7,-17380.,-186.82,-20904.,-6472.6,-4539.4,-3033.4,67.465,2403.4,2191.5,1416.6,333.93,2992.6,1686.6,0.0000,6616.9,4449.7,4252.8,3658.0,0.0000,-402.29,-127.77,-83.158,-45.009,-116.59,-587.69,0.0000,-1084.7,-1628.6,-759.17,-1329.8
519.0000000000,97.549,2005.6,2084.6,1362.1,304.33,2788.4,973.62,0.91901,5508.2,2621.8,3350.5,1945.3,0.0000,-8021.9,-7416.1,-1805.7,-2804.7,-3491.2,-17376.,-186.57,-20897.,-6472.3,-4538.7,-3032.4,67.286,2397.0,2185.7,1410.5,333.00,2978.8,1686.6,0.0000,6608.5,4449.7,4252.8,3658.0,0.0000,-401.06,-127.37,-82.858,-44.885,-115.89,-587.69,0.0000,-1084.5,-1628.3,-759.16,-1329.5
520.0000000000,97.366,2001.7,2080.3,1357.3,303.54,2779.6,973.62,0.91958,5503.0,2622.0,3350.6,1945.6,0.0000,-8014.8,-7413.8,-1802.8,-2802.8,-3483.8,-17372.,-186.33,-20890.,-6472.0,-4538.1,-3031.4,67.104,2390.5,2179.8,1404.4,332.06,2965.0,1686.6,0.0000,6600.2,4449.7,4252.8,3658.0,0.0000,-399.80,-126.95,-82.555,-44.758,-115.20,-587.69,0.0000,-1084.4,-1628.1,-759.14,-1329.2
521.0000000000,97.178,1997.2,2075.4,1352.6,302.73,2768.5,973.62,0.92012,5496.5,2622.2,3350.6,1945.9,0.0000,-8007.4,-7411.3,-1799.8,-2801.0,-3476.3,-17368.,-186.08,-20884.,-6471.7,-4537.4,-3030.4,66.909,2383.6,2173.5,1398.2,331.06,2951.1,1686.6,0.0000,6591.7,4449.7,4252.8,3658.0,0.0000,-398.46,-126.51,-82.243,-44.623,-114.50,-587.69,0.0000,-1084.2,-1627.9,-759.13,-1328.9
522.0000000000,96.980,1993.4,2070.6,1347.2,301.88,2756.4,973.62,0.92068,5489.4,2622.4,3350.6,1946.2,0.0000,-7999.9,-7408.8,-1796.9,-2799.1,-3468.8,-17365.,-185.84,-20877.,-6471.4,-4536.7,-3029.4,66.714,2376.7,2167.1,1392.1,330.06,2937.3,1686.6,0.0000,6583.4,4449.7,4252.8,3658.0,0.0000,-397.13,-126.06,-81.932,-44.487,-113.81,-587.69,0.0000,-1084.1,-1627.7,-759.12,-1328.6
523.0000000000,96.780,1988.6,2066.0,1341.6,301.03,2743.7,973.62,0.93207,5481.6,2622.7,3350.6,1946.4,0.0000,-7992.2,-7406.2,-1793.9,-2797.2,-3461.4,-17361.,-185.59,-20870.,-6471.1,-4536.1,-3028.4,66.520,2369.7,2160.8,1386.0,329.06,2923.7,1686.6,0.0000,6575.1,4449.7,4252.8,3658.0,0.0000,-395.79,-125.62,-81.624,-44.352,-113.13,-587.69,0.0000,-1083.9,-1627.5,-759.11,-1328.3
524.0000000000,96.577,1983.6,2060.9,1335.9,300.15,2731.2,973.62,0.93612,5473.8,2622.9,3350.6,1946.7,0.0000,-7984.3,-7403.6,-1791.0,-2795.3,-3453.9,-17357.,-185.35,-20864.,-6470.8,-4535.4,-3027.4,66.329,2362.9,2154.6,1380.0,328.09,2910.3,1686.6,0.0000,6567.1,4449.7,4252.8,3658.0,0.0000,-394.47,-125.19,-81.321,-44.219,-112.46,-587.69,0.0000,-1083.8,-1627.2,-759.10,-1328.1
525.0000000000,96.529,1978.8,2055.8,1330.1,299.31,2719.3,973.62,0.93668,5466.4,2623.1,3350.6,1947.0,0.0000,-7976.4,-7401.0,-1788.0,-2793.4,-3446.4,-17353.,-185.11,-20857.,-6470.5,-4534.8,-3026.4,66.162,2357.0,2149.2,1374.6,327.23,2898.1,1686.6,0.0000,6559.7,4449.7,4252.8,3658.0,0.0000,-393.30,-124.79,-81.049,-44.108,-111.83,-587.69,0.0000,-1083.6,-1627.0,-759.08,-1327.8
526.0000000000,96.379,1974.1,2051.1,1324.6,298.54,2707.7,973.62,0.93724,5459.3,2623.3,3350.6,1947.3,0.0000,-7968.5,-7398.3,-1785.0,-2791.5,-3438.9,-17349.,-184.86,-20850.,-6470.2,-4534.1,-3025.4,66.016,2351.8,2144.5,1369.3,326.47,2886.1,1686.6,0.0000,6552.4,4449.7,4252.8,3658.0,0.0000,-392.25,-124.44,-80.795,-44.011,-111.21,-587.69,0.0000,-1083.5,-1626.8,-759.07,-1327.5
527.0000000000,96.204,1970.0,2046.2,1319.3,297.79,2696.7,973.62,0.93776,5451.9,2623.5,3350.6,1947.6,0.0000,-7960.5,-7395.5,-1782.0,-2789.6,-3431.4,-17345.,-184.62,-20843.,-6469.9,-4533.4,-3024.4,65.832,2345.2,2138.4,1363.5,325.52,2873.1,1686.6,0.0000,6544.6,4449.7,4252.8,3658.0,0.0000,-390.98,-124.02,-80.502,-43.888,-110.56,-587.69,0.0000,-1083.4,-1626.6,-759.06,-1327.2
528.0000000000,96.018,1965.4,2041.1,1313.8,297.03,2685.1,973.62,0.94377,5444.4,2623.8,3350.6,1947.9,0.0000,-7952.4,-7392.8,-1779.0,-2787.7,-3424.0,-17341.,-184.38,-20836.,-6469.6,-4532.7,-3023.4,65.672,2339.5,2133.3,1358.1,324.70,2861.0,1686.6,0.0000,6537.2,4449.7,4252.8,3658.0,0.0000,-389.87,-123.64,-80.236,-43.781,-109.94,-587.69,0.0000,-1083.2,-1626.4,-759.04,-1326.9
529.0000000000,95.847,1960.5,2035.7,1308.7,296.30,2673.4,973.59,0.95443,5437.3,2624.0,3350.7,1948.2,0.0000,-7944.3,-7390.0,-1776.0,-2785.8,-3416.5,-17337.,-184.14,-20830.,-6469.2,-4532.1,-3022.4,65.495,2333.2,2127.5,1352.9,323.80,2849.4,1686.6,10.304,6530.4,4452.2,4252.8,3658.9,0.0000,-388.66,-123.22,-79.966,-43.663,-109.34,-587.69,-0.47191,-1083.1,-1626.2,-759.03,-1326.7
530.0000000000,95.679,1958.6,2033.5,1303.8,296.08,2662.0,973.53,0.95499,5430.4,2624.2,3350.7,1948.4,0.0000,-7936.3,-7387.3,-1773.1,-2783.9,-3409.1,-17334.,-183.90,-20823.,-6468.9,-4531.4,-3021.4,73.926,2357.7,2149.5,1357.2,327.51,2852.3,1686.6,0.0000,6532.0,4449.7,4252.8,3658.0,0.0000,-391.51,-124.22,-80.330,-44.009,-109.29,-587.69,0.0000,-1083.1,-1625.9,-759.02,-1326.4
531.0000000000,95.855,1962.5,2035.7,1299.6,296.70,2652.4,973.53,0.95556,5423.7,2624.4,3350.7,1948.7,0.0000,-7928.9,-7384.9,-1770.2,-2782.1,-3401.7,-17330.,-183.66,-20816.,-6468.5,-4530.7,-3020.4,66.007,2351.5,2144.1,1351.4,326.12,2839.7,1686.6,0.0000,6524.2,4449.7,4252.8,3658.0,0.0000,-391.38,-124.04,-80.177,-44.005,-108.67,-587.69,0.0000,-1082.9,-1625.7,-759.01,-1326.1
532.0000000000,95.855,1963.9,2037.0,1296.6,296.70,2643.3,973.53,0.95612,5417.5,2624.6,3350.6,1949.0,0.0000,-7921.8,-7382.6,-1767.3,-2780.4,-3394.4,-17326.,-183.43,-20809.,-6468.2,-4530.0,-3019.4,65.920,2348.4,2141.3,1346.2,325.63,2827.1,1686.6,0.0000,6516.5,4449.7,4252.8,3658.0,0.0000,-390.71,-123.81,-79.953,-43.947,-108.03,-587.69,0.0000,-1082.8,-1625.5,-758.99,-1325.8
533.0000000000,95.869,1962.6,2035.8,1293.2,296.86,2633.4,973.53,0.95666,5411.1,2624.9,3350.6,1949.3,0.0000,-7914.7,-7380.4,-1764.5,-2778.6,-3387.1,-17322.,-183.19,-20803.,-6467.8,-4529.3,-3018.4,65.799,2344.1,2137.4,1340.9,324.98,2814.6,1686.6,0.0000,6509.0,4449.7,4252.8,3658.0,0.0000,-389.84,-123.51,-79.709,-43.866,-107.40,-587.69,0.0000,-1082.6,-1625.3,-758.98,-1325.5
534.0000000000,95.856,1959.9,2033.8,1289.1,296.42,2623.5,973.53,0.95721,5404.7,2625.1,3350.6,1949.6,0.0000,-7907.6,-7378.0,-1761.6,-2776.8,-3379.8,-17318.,-182.95,-20796.,-6467.4,-4528.6,-3017.3,65.655,2338.9,2132.7,1335.4,324.23,2802.2,1686.6,0.0000,6501.4,4449.7,4252.8,3658.0,0.0000,-388.84,-123.17,-79.449,-43.770,-106.78,-587.69,0.0000,-1082.5,-1625.1,-758.97,-1325.3
535.0000000000,95.739,1956.9,2031.3,1284.6,295.82,2613.0,973.53,0.95775,5398.7,2625.3,3350.6,1949.8,0.0000,-7900.4,-7375.6,-1758.7,-2775.0,-3372.4,-17314.,-182.71,-20789.,-6467.1,-4528.0,-3016.3,65.505,2333.6,2127.8,1330.1,323.45,2790.0,1686.6,0.0000,6494.1,4449.7,4252.8,3658.0,0.0000,-387.80,-122.82,-79.190,-43.670,-106.16,-587.69,0.0000,-1082.4,-1624.9,-758.95,-1325.0
536.0000000000,95.694,1968.6,2042.2,1281.1,297.92,2605.3,973.53,0.95832,5393.2,2625.5,3350.6,1950.1,0.0000,-7894.4,-7373.8,-1756.1,-2773.3,-3365.2,-17310.,-182.48,-20783.,-6466.7,-4527.3,-3015.4,135.52,2511.8,2285.0,1382.3,343.16,2882.2,1686.8,236.59,6550.2,4457.6,4254.3,3661.2,0.0000,-405.99,-129.75,-82.401,-45.750,-109.51,-587.69,-10.836,-1082.9,-1624.7,-758.95,-1324.9
537.0000000000,97.327,2016.2,2083.1,1291.7,305.48,2628.8,973.53,0.95890,5394.0,2625.7,3350.6,1950.4,0.0000,-7892.3,-7374.1,-1754.9,-2772.0,-3359.0,-17307.,-182.26,-20777.,-6466.4,-4526.6,-3014.4,761.94,3171.9,3130.7,1652.8,381.64,3518.6,1691.1,383.44,6954.5,4580.8,4313.1,3756.8,0.0000,-422.35,-150.86,-92.104,-47.630,-133.35,-587.76,-17.562,-1087.4,-1624.4,-759.24,-1329.7
538.0000000000,99.078,2070.8,2136.3,1342.3,314.12,2720.5,973.53,0.95947,5413.5,2625.9,3350.6,1950.6,0.0000,-7893.9,-7376.5,-1756.0,-2771.1,-3355.4,-17303.,-182.04,-20773.,-6466.0,-4525.9,-3013.4,72.630,2587.4,2359.3,1712.8,444.59,3717.7,1708.7,134.17,7103.2,4667.3,4484.7,3897.2,0.0000,-429.72,-136.12,-94.474,-48.948,-137.97,-588.06,-6.1452,-1089.3,-1624.2,-760.12,-1336.8
539.0000000000,100.74,2108.1,2174.3,1413.6,324.45,2829.5,973.53,0.96002,5444.4,2626.1,3350.9,1950.9,0.0000,-7897.2,-7379.6,-1757.8,-2770.3,-3355.5,-17299.,-181.82,-20771.,-6465.7,-4525.2,-3012.4,72.800,2593.4,2364.8,1695.6,379.14,3646.2,1686.6,0.0000,7025.4,4470.5,4272.2,3666.0,0.0000,-430.70,-136.47,-95.042,-48.636,-138.65,-587.69,0.0000,-1088.0,-1624.0,-759.00,-1324.3
540.0000000000,101.89,2124.8,2194.1,1469.6,328.30,2910.2,973.53,0.96056,5475.0,2626.3,3350.8,1951.3,0.0000,-7900.4,-7382.4,-1760.7,-2769.4,-3357.8,-17295.,-181.58,-20769.,-6465.3,-4524.5,-3011.4,72.765,2592.2,2363.7,1697.9,366.83,3661.7,1686.6,0.0000,7026.0,4454.5,4257.3,3659.0,0.0000,-430.47,-136.42,-95.423,-48.534,-139.71,-587.69,0.0000,-1087.9,-1623.8,-758.91,-1323.7
541.0000000000,102.53,2139.3,2209.6,1521.7,330.80,2970.8,973.53,0.96111,5494.8,2626.6,3350.7,1951.7,0.0000,-7903.4,-7384.9,-1763.5,-2768.5,-3358.8,-17291.,-181.36,-20767.,-6464.9,-4523.8,-3010.4,537.14,3208.3,2975.5,1839.8,502.84,3899.5,1719.3,510.99,7229.7,4671.5,4464.2,3888.2,0.0000,-438.72,-150.95,-97.410,-50.176,-144.02,-588.23,-23.404,-1090.6,-1623.6,-759.98,-1335.5
542.0000000000,103.34,2161.1,2230.2,1556.8,333.74,3026.0,973.51,0.96166,5528.2,2626.8,3351.2,1952.6,0.0000,-7907.0,-7387.7,-1767.5,-2767.6,-3359.1,-17287.,-181.13,-20765.,-6464.6,-4523.1,-3009.5,74.410,2650.8,2417.1,1766.1,385.81,3815.0,1686.6,0.0000,7120.4,4451.5,4255.9,3658.3,0.0000,-440.22,-139.58,-98.239,-49.698,-144.90,-587.69,0.0000,-1088.9,-1623.4,-758.88,-1323.1
543.0000000000,103.67,2175.1,2248.0,1594.2,335.69,3069.9,973.50,0.96222,5568.0,2627.0,3351.8,1954.1,0.0000,-7910.7,-7390.5,-1771.8,-2766.7,-3359.1,-17284.,-180.89,-20764.,-6464.2,-4522.4,-3008.5,74.395,2650.3,2416.6,1766.2,372.20,3822.7,1686.6,0.0000,7120.4,4449.7,4252.9,3658.0,0.0000,-440.15,-139.60,-98.675,-49.600,-146.05,-587.69,0.0000,-1088.7,-1623.2,-758.85,-1322.9
544.0000000000,104.02,2183.3,2258.4,1614.1,336.94,3142.4,973.46,0.96275,5650.6,2628.4,3351.3,1953.8,0.0000,-7914.2,-7392.9,-1775.1,-2765.7,-3358.9,-17280.,-180.66,-20763.,-6463.9,-4521.6,-3007.5,74.256,2645.3,2412.1,1776.8,371.27,3851.7,1686.6,0.0000,7137.9,4449.7,4252.8,3658.0,0.0000,-439.35,-139.37,-98.980,-49.504,-147.21,-587.69,0.0000,-1088.9,-1623.0,-758.83,-1322.6
545.0000000000,104.09,2185.5,2262.4,1630.6,336.99,3236.8,973.45,0.96326,5721.0,2629.3,3351.6,1954.1,0.0000,-7917.1,-7394.8,-1777.7,-2764.6,-3358.4,-17276.,-180.43,-20762.,-6463.5,-4520.9,-3006.5,74.055,2638.2,2405.6,1786.1,370.50,3878.2,1686.6,0.0000,7154.0,4449.7,4252.8,3658.0,0.0000,-438.17,-139.03,-99.195,-49.370,-148.24,-587.69,0.0000,-1089.0,-1622.8,-758.82,-1322.3
546.0000000000,103.71,2184.2,2260.2,1648.0,336.49,3312.3,973.43,0.96380,5770.4,2629.4,3351.8,1954.3,0.0000,-7919.0,-7396.3,-1780.1,-2763.5,-3357.8,-17273.,-180.19,-20760.,-6463.2,-4520.2,-3005.5,73.819,2629.8,2397.9,1794.0,369.56,3901.5,1686.6,0.0000,7168.2,4449.7,4252.8,3658.0,0.0000,-436.78,-138.61,-99.346,-49.213,-149.14,-587.69,0.0000,-1089.1,-1622.6,-758.80,-1322.1
547.0000000000,103.51,2183.3,2256.8,1666.0,335.80,3353.3,973.39,0.96433,5805.5,2629.8,3351.8,1954.3,0.0000,-7920.0,-7397.4,-1782.3,-2762.3,-3357.1,-17269.,-179.96,-20759.,-6462.8,-4519.5,-3004.5,73.585,2621.4,2390.3,1801.2,368.60,3922.8,1686.6,0.0000,7181.3,4449.7,4252.8,3658.0,0.0000,-435.39,-138.18,-99.473,-49.057,-149.97,-587.69,0.0000,-1089.2,-1622.4,-758.79,-1321.8
548.0000000000,103.44,2180.5,2255.0,1678.2,335.00,3387.2,973.35,0.96485,5834.3,2629.9,3352.6,1954.7,0.0000,-7920.2,-7398.2,-1784.2,-2761.1,-3356.4,-17265.,-179.73,-20758.,-6462.5,-4518.8,-3003.5,73.340,2612.7,2382.3,1807.4,367.59,3941.6,1686.6,0.0000,7192.8,4449.7,4252.8,3658.0,0.0000,-433.92,-137.74,-99.559,-48.893,-150.70,-587.69,0.0000,-1089.2,-1622.2,-758.78,-1321.6
549.0000000000,103.30,2176.3,2251.1,1688.3,334.16,3411.9,973.35,0.96537,5852.9,2629.9,3352.6,1954.7,0.0000,-7919.8,-7398.7,-1785.9,-2759.8,-3355.7,-17262.,-179.50,-20757.,-6462.2,-4518.1,-3002.5,73.093,2603.9,2374.3,1812.8,366.54,3958.6,1686.6,0.0000,7203.1,4449.7,4252.8,3658.0,0.0000,-432.44,-137.28,-99.618,-48.728,-151.35,-587.69,0.0000,-1089.3,-1622.0,-758.76,-1321.3
550.0000000000,103.16,2171.6,2246.1,1696.1,333.29,3434.4,973.35,0.96587,5866.9,2631.3,3352.1,1955.0,0.0000,-7918.9,-7398.9,-1787.4,-2758.5,-3355.0,-17258.,-179.26,-20757.,-6461.9,-4517.4,-3001.5,72.841,2594.9,2366.1,1817.2,365.46,3972.8,1686.6,0.0000,7211.8,4449.7,4252.8,3658.0,0.0000,-430.92,-136.80,-99.639,-48.561,-151.90,-587.69,0.0000,-1089.3,-1621.8,-758.75,-1321.0
551.0000000000,102.90,2166.4,2242.4,1702.5,332.39,3466.0,973.31,0.96641,5887.0,2632.0,3351.7,1955.2,0.0000,-7917.6,-7398.9,-1788.8,-2757.2,-3354.4,-17255.,-179.03,-20756.,-6461.6,-4516.7,-3000.5,72.585,2585.8,2357.8,1820.7,364.35,3984.8,1686.6,0.0000,7219.2,4449.7,4252.8,3658.0,0.0000,-429.37,-136.32,-99.628,-48.390,-152.37,-587.69,0.0000,-1089.4,-1621.6,-758.74,-1320.8
552.0000000000,102.64,2161.6,2236.9,1710.2,331.47,3489.4,973.30,0.96693,5905.7,2632.3,3351.7,1955.3,0.0000,-7915.8,-7398.7,-1790.1,-2755.8,-3354.0,-17251.,-178.80,-20755.,-6461.3,-4516.0,-2999.5,72.330,2576.7,2349.5,1823.5,363.23,3994.8,1686.6,0.0000,7225.3,4449.7,4252.8,3658.0,0.0000,-427.81,-135.83,-99.591,-48.220,-152.75,-587.69,0.0000,-1089.4,-1621.4,-758.73,-1320.5
553.0000000000,102.38,2155.6,2230.2,1717.3,330.52,3514.2,973.29,0.96744,5915.6,2631.9,3351.6,1955.7,0.0000,-7913.4,-7398.2,-1791.2,-2754.4,-3353.6,-17248.,-178.57,-20753.,-6461.0,-4515.3,-2998.5,72.071,2567.5,2341.1,1825.4,362.07,4002.7,1686.6,0.0000,7230.2,4449.7,4252.8,3658.0,0.0000,-426.22,-135.32,-99.523,-48.047,-153.05,-587.69,0.0000,-1089.4,-1621.2,-758.71,-1320.3
554.0000000000,102.11,2149.0,2223.8,1721.5,329.54,3532.4,973.29,0.96796,5924.8,2630.9,3351.6,1955.8,0.0000,-7910.7,-7397.5,-1792.2,-2753.0,-3353.2,-17244.,-178.34,-20752.,-6460.7,-4514.6,-2997.5,71.812,2558.3,2332.7,1826.6,360.90,4008.8,1686.6,0.0000,7233.9,4449.7,4252.8,3658.0,0.0000,-424.63,-134.82,-99.432,-47.875,-153.28,-587.69,0.0000,-1089.4,-1621.0,-758.70,-1320.0
555.0000000000,101.84,2141.9,2217.0,1725.1,328.56,3544.1,973.29,0.96847,5938.6,2631.0,3351.9,1955.9,0.0000,-7907.6,-7396.6,-1793.1,-2751.6,-3352.8,-17241.,-178.11,-20751.,-6460.4,-4513.9,-2996.5,71.555,2549.1,2324.4,1827.2,359.73,4013.2,1686.6,0.0000,7236.7,4449.7,4252.8,3658.0,0.0000,-423.04,-134.31,-99.320,-47.704,-153.44,-587.69,0.0000,-1089.3,-1620.8,-758.69,-1319.8
556.0000000000,101.58,2135.5,2209.8,1727.3,327.58,3553.2,973.29,0.96898,5949.7,2631.2,3351.9,1956.0,0.0000,-7904.1,-7395.5,-1793.8,-2750.1,-3352.2,-17237.,-177.88,-20750.,-6460.1,-4513.2,-2995.5,71.317,2540.6,2316.6,1827.3,358.64,4016.4,1686.6,0.0000,7238.6,4449.7,4252.8,3658.0,0.0000,-421.56,-133.83,-99.204,-47.545,-153.55,-587.69,0.0000,-1089.3,-1620.6,-758.67,-1319.5
557.0000000000,101.32,2129.5,2202.8,1729.3,326.63,3567.4,973.29,0.96948,5958.9,2631.4,3351.9,1956.5,0.0000,-7900.2,-7394.2,-1794.4,-2748.6,-3351.8,-17234.,-177.65,-20749.,-6459.8,-4512.5,-2994.5,71.084,2532.3,2309.1,1827.3,357.57,4018.8,1686.6,0.0000,7240.1,4449.7,4252.8,3658.0,0.0000,-420.10,-133.36,-99.082,-47.389,-153.63,-587.69,0.0000,-1089.3,-1620.4,-758.66,-1319.2
558.0000000000,101.08,2124.1,2198.0,1731.3,325.92,3574.9,973.29,0.96999,5967.8,2631.6,3351.8,1956.8,0.0000,-7896.2,-7392.7,-1795.0,-2747.1,-3351.4,-17231.,-177.42,-20747.,-6459.4,-4511.8,-2993.5,71.096,2537.7,2309.4,1830.3,357.68,4026.6,1686.6,0.0000,7244.9,4449.7,4252.8,3658.0,0.0000,-420.10,-133.34,-99.192,-47.397,-153.92,-587.69,0.0000,-1089.3,-1620.2,-758.65,-1319.0
559.0000000000,100.96,2120.2,2195.1,1732.5,325.41,3585.5,973.29,0.89930,5973.6,2631.8,3351.7,1957.0,0.0000,-7892.1,-7391.3,-1795.4,-2745.6,-3351.0,-17227.,-177.19,-20746.,-6459.1,-4511.1,-2992.6,70.850,2524.0,2301.5,1828.8,356.52,4025.3,1686.6,0.0000,7244.2,4449.7,4252.8,3658.0,0.0000,-418.55,-132.84,-99.013,-47.234,-153.85,-587.69,0.0000,-1089.2,-1620.0,-758.64,-1318.7
560.0000000000,100.90,2115.3,2192.9,1733.2,324.62,3596.8,973.29,0.77122,5980.8,2632.0,3351.7,1957.2,0.0000,-7888.0,-7389.6,-1795.7,-2744.2,-3350.5,-17224.,-176.97,-20744.,-6458.8,-4510.4,-2991.6,70.600,2515.1,2293.4,1826.6,355.34,4022.6,1686.6,0.0000,7242.5,4449.7,4252.8,3658.0,0.0000,-416.98,-132.33,-98.811,-47.067,-153.73,-587.69,0.0000,-1089.2,-1619.8,-758.62,-1318.5
561.0000000000,100.74,2109.1,2186.5,1733.3,323.83,3600.3,973.29,2.5070,5996.8,2632.2,3351.7,1957.4,0.0000,-7883.6,-7387.8,-1796.0,-2742.6,-3349.8,-17221.,-176.74,-20743.,-6458.4,-4509.7,-2990.6,70.350,2506.2,2285.2,1824.0,354.15,4018.6,1686.6,0.0000,7240.1,4449.7,4252.8,3658.0,0.0000,-415.41,-131.82,-98.592,-46.900,-153.55,-587.69,0.0000,-1089.1,-1619.6,-758.61,-1318.2
562.0000000000,100.51,2102.4,2179.9,1733.0,322.84,3604.4,973.29,2.5244,6002.7,2632.3,3351.5,1957.5,0.0000,-7879.0,-7385.9,-1796.1,-2741.1,-3349.0,-17218.,-176.51,-20741.,-6458.1,-4509.0,-2989.6,70.132,2498.4,2278.1,1823.3,353.13,4019.1,1686.6,189.14,7258.4,4507.7,4278.6,3728.6,0.0000,-414.02,-131.36,-98.455,-46.754,-153.55,-587.69,-8.6629,-1089.3,-1619.4,-758.73,-1321.5
563.0000000000,100.28,2097.8,2177.8,1732.8,322.24,3611.9,973.26,2.5247,6007.8,2632.3,3351.3,1957.9,0.0000,-7874.4,-7383.9,-1796.2,-2739.6,-3348.0,-17214.,-176.29,-20739.,-6457.8,-4508.3,-2988.6,75.603,2519.7,2295.0,1831.9,358.06,4034.1,1686.6,0.0000,7250.9,4449.7,4252.8,3658.0,0.0000,-414.79,-131.84,-98.688,-46.876,-153.96,-587.69,0.0000,-1089.1,-1619.2,-758.58,-1317.7
564.0000000000,100.24,2097.4,2178.3,1732.9,322.28,3617.7,973.25,2.5251,6014.5,2632.5,3351.3,1958.1,0.0000,-7870.1,-7382.0,-1796.2,-2738.0,-3347.2,-17211.,-176.07,-20737.,-6457.4,-4507.6,-2987.6,73.627,2506.5,2295.4,1830.5,362.03,4035.3,1686.6,0.0000,7250.3,4449.7,4252.8,3658.0,0.0000,-415.16,-131.90,-98.819,-46.955,-154.14,-587.69,0.0000,-1089.1,-1619.0,-758.57,-1317.4
565.0000000000,100.21,2096.7,2177.4,1733.8,322.22,3626.1,973.23,2.5254,6017.4,2632.7,3351.4,1958.2,0.0000,-7866.0,-7380.3,-1796.3,-2736.6,-3346.8,-17208.,-175.84,-20736.,-6457.1,-4506.9,-2986.7,70.183,2500.2,2279.8,1826.9,353.43,4028.0,1686.6,0.0000,7245.9,4449.7,4252.8,3658.0,0.0000,-414.03,-131.32,-98.606,-46.789,-153.82,-587.69,0.0000,-1089.0,-1618.8,-758.55,-1317.2
566.0000000000,100.12,2093.2,2174.1,1734.2,321.89,3631.9,973.20,2.5258,6018.7,2632.9,3351.4,1958.5,0.0000,-7861.7,-7378.5,-1796.2,-2735.1,-3346.2,-17205.,-175.62,-20734.,-6456.7,-4506.2,-2985.8,69.977,2492.9,2273.1,1822.6,352.41,4019.1,1686.6,0.0000,7240.5,4449.7,4252.8,3658.0,0.0000,-412.71,-130.88,-98.352,-46.651,-153.45,-587.69,0.0000,-1088.9,-1618.6,-758.54,-1316.9
567.0000000000,100.01,2088.2,2169.4,1732.9,321.25,3632.3,973.20,2.5324,6019.0,2633.0,3351.4,1958.8,0.0000,-7857.2,-7376.5,-1796.1,-2733.5,-3345.3,-17202.,-175.40,-20732.,-6456.4,-4505.5,-2984.9,69.756,2485.0,2265.9,1817.8,351.31,4009.2,1686.6,0.0000,7234.5,4449.7,4252.8,3658.0,0.0000,-411.30,-130.42,-98.075,-46.504,-153.04,-587.69,0.0000,-1088.8,-1618.4,-758.53,-1316.6
568.0000000000,99.823,2082.5,2163.7,1730.3,320.35,3630.9,973.20,2.5424,6019.0,2633.1,3351.4,1959.1,0.0000,-7852.4,-7374.4,-1795.8,-2732.0,-3344.1,-17199.,-175.17,-20730.,-6456.0,-4504.8,-2983.9,69.528,2476.9,2258.5,1812.7,350.18,3998.4,1686.6,0.0000,7228.1,4449.7,4252.8,3658.0,0.0000,-409.85,-129.94,-97.783,-46.352,-152.59,-587.69,0.0000,-1088.7,-1618.2,-758.51,-1316.4
569.0000000000,99.596,2076.6,2157.7,1726.7,319.41,3632.1,973.20,1.2488,6019.3,2633.4,3351.4,1959.3,0.0000,-7847.4,-7372.1,-1795.4,-2730.4,-3342.7,-17195.,-174.95,-20727.,-6455.7,-4504.1,-2983.0,69.304,2468.9,2251.2,1807.4,349.06,3987.2,1686.6,0.0000,7221.3,4449.7,4252.8,3658.0,0.0000,-408.42,-129.47,-97.486,-46.203,-152.12,-587.69,0.0000,-1088.5,-1618.0,-758.50,-1316.1
570.0000000000,99.361,2070.3,2151.8,1722.3,318.44,3629.3,973.20,0.95801,6019.0,2633.8,3351.2,1959.5,0.0000,-7842.0,-7369.8,-1794.9,-2728.8,-3341.1,-17192.,-174.72,-20725.,-6455.3,-4503.4,-2982.0,69.077,2460.8,2243.9,1801.8,347.92,3975.2,1686.6,0.0000,7214.0,4449.7,4252.8,3658.0,0.0000,-406.97,-128.99,-97.177,-46.051,-151.61,-587.69,0.0000,-1088.4,-1617.8,-758.48,-1315.9
571.0000000000,99.115,2064.8,2146.2,1717.9,317.58,3628.7,973.20,0.95849,6017.8,2634.0,3351.2,1959.7,0.0000,-7836.6,-7367.4,-1794.3,-2727.2,-3339.4,-17189.,-174.50,-20723.,-6454.9,-4502.7,-2981.1,68.989,2457.7,2241.0,1798.4,347.46,3967.3,1686.6,0.0000,7209.3,4449.7,4252.8,3658.0,0.0000,-406.34,-128.77,-97.016,-45.993,-151.27,-587.69,0.0000,-1088.3,-1617.6,-758.47,-1315.6
572.0000000000,98.953,2060.3,2140.7,1713.8,316.84,3624.7,973.12,0.95897,6019.8,2634.2,3351.2,1960.0,0.0000,-7831.0,-7365.0,-1793.6,-2725.7,-3337.4,-17186.,-174.28,-20721.,-6454.6,-4502.0,-2980.1,68.763,2449.7,2233.7,1792.3,346.32,3954.2,1686.6,0.0000,7201.3,4449.7,4252.8,3658.0,0.0000,-404.89,-128.29,-96.693,-45.842,-150.72,-587.69,0.0000,-1088.2,-1617.4,-758.45,-1315.4
573.0000000000,98.733,2054.8,2134.8,1709.4,315.94,3618.8,973.12,1.0261,6016.1,2634.2,3351.2,1960.2,0.0000,-7825.3,-7362.6,-1792.8,-2724.0,-3335.4,-17183.,-174.06,-20719.,-6454.2,-4501.3,-2979.2,68.533,2441.4,2226.2,1786.0,345.15,3940.3,1686.6,0.0000,7192.9,4449.7,4252.8,3658.0,0.0000,-403.41,-127.80,-96.358,-45.689,-150.13,-587.69,0.0000,-1088.1,-1617.2,-758.44,-1315.2
574.0000000000,98.526,2048.9,2128.1,1704.5,315.04,3614.7,973.12,2.7136,6014.3,2634.4,3351.2,1960.5,0.0000,-7819.3,-7360.0,-1791.9,-2722.4,-3333.2,-17180.,-173.84,-20717.,-6453.8,-4500.6,-2978.2,68.302,2433.2,2218.7,1779.4,343.99,3925.9,1686.6,0.0000,7184.2,4449.7,4252.8,3658.0,0.0000,-401.93,-127.31,-96.015,-45.535,-149.52,-587.69,0.0000,-1087.9,-1617.0,-758.43,-1314.9
575.0000000000,98.303,2042.7,2121.7,1699.1,314.04,3605.9,973.06,2.4677,6009.6,2634.3,3351.3,1960.8,0.0000,-7813.1,-7357.4,-1790.9,-2720.8,-3330.8,-17177.,-173.62,-20715.,-6453.5,-4499.9,-2977.2,68.079,2425.3,2211.4,1772.9,342.85,3911.3,1686.6,0.0000,7175.4,4449.7,4252.8,3658.0,0.0000,-400.49,-126.83,-95.675,-45.386,-148.91,-587.69,0.0000,-1087.8,-1616.8,-758.41,-1314.7
576.0000000000,98.068,2036.4,2115.0,1693.5,313.06,3596.3,973.03,1.1285,6004.4,2634.7,3351.2,1961.0,0.0000,-7806.8,-7354.8,-1789.9,-2719.2,-3328.3,-17174.,-173.40,-20712.,-6453.1,-4499.2,-2976.3,67.854,2417.2,2204.1,1766.0,341.70,3896.2,1686.6,0.0000,7166.2,4449.7,4252.8,3658.0,0.0000,-399.04,-126.34,-95.326,-45.236,-148.26,-587.69,0.0000,-1087.7,-1616.6,-758.40,-1314.4
577.0000000000,97.832,2030.2,2108.6,1687.5,312.06,3586.3,973.03,1.1291,6001.9,2635.0,3351.3,1961.3,0.0000,-7800.2,-7352.0,-1788.7,-2717.5,-3325.6,-17170.,-173.18,-20709.,-6452.7,-4498.5,-2975.3,67.629,2409.2,2196.8,1759.1,340.54,3880.6,1686.6,0.0000,7156.8,4449.7,4252.8,3658.0,0.0000,-397.59,-125.86,-94.972,-45.086,-147.60,-587.69,0.0000,-1087.5,-1616.4,-758.38,-1314.2
578.0000000000,97.598,2023.9,2102.1,1681.3,311.07,3575.4,973.03,1.1297,5999.4,2635.2,3351.3,1961.6,0.0000,-7793.6,-7349.3,-1787.5,-2715.9,-3322.9,-17167.,-172.96,-20707.,-6452.3,-4497.8,-2974.3,67.414,2401.6,2189.8,1752.1,339.44,3865.0,1686.6,0.0000,7147.4,4449.7,4252.8,3658.0,0.0000,-396.19,-125.39,-94.624,-44.942,-146.94,-587.69,0.0000,-1087.4,-1616.2,-758.37,-1313.9
579.0000000000,97.371,2018.3,2096.0,1675.2,310.17,3564.3,973.01,1.1303,5996.2,2635.5,3351.3,1961.8,0.0000,-7786.9,-7346.5,-1786.2,-2714.2,-3320.0,-17164.,-172.75,-20704.,-6452.0,-4497.1,-2973.4,67.285,2397.0,2185.7,1749.8,338.80,3859.4,1686.6,100.57,7151.1,4461.7,4260.6,3671.2,0.0000,-395.30,-125.09,-94.465,-44.857,-146.66,-587.69,-4.6060,-1087.4,-1616.0,-758.39,-1314.3
580.0000000000,97.231,2020.8,2097.1,1670.9,310.76,3556.6,973.00,1.1308,5990.7,2635.9,3351.3,1962.1,0.0000,-7780.8,-7344.0,-1785.1,-2712.6,-3317.1,-17161.,-172.54,-20701.,-6451.6,-4496.4,-2972.4,80.199,2465.7,2249.4,1777.5,350.55,3909.7,1686.6,652.16,7198.3,4486.4,4279.5,3696.7,0.0000,-403.31,-127.99,-95.984,-45.807,-148.41,-587.69,-29.870,-1087.9,-1615.8,-758.48,-1315.3
581.0000000000,97.873,2037.7,2110.0,1671.3,313.41,3555.9,973.00,1.1314,5986.8,2636.1,3351.3,1962.3,0.0000,-7776.2,-7342.4,-1784.2,-2711.2,-3314.4,-17158.,-172.33,-20698.,-6451.2,-4495.7,-2971.5,69.068,2460.5,2243.6,1770.8,347.48,3894.6,1686.6,0.0000,7166.2,4454.7,4252.8,3658.4,0.0000,-405.55,-128.30,-96.109,-46.046,-147.90,-587.69,0.0000,-1087.5,-1615.6,-758.32,-1313.2
582.0000000000,98.187,2049.0,2121.4,1675.8,314.80,3554.5,973.00,1.1352,5983.5,2636.2,3351.4,1962.6,0.0000,-7772.4,-7341.3,-1783.3,-2709.8,-3312.0,-17155.,-172.12,-20695.,-6450.9,-4495.0,-2970.5,69.070,2460.6,2243.6,1764.6,347.28,3878.6,1686.6,0.0000,7155.3,4450.1,4252.8,3658.0,0.0000,-405.46,-128.26,-95.899,-46.047,-147.22,-587.69,0.0000,-1087.3,-1615.4,-758.31,-1312.9
583.0000000000,98.503,2052.6,2124.8,1677.2,316.07,3548.5,973.00,1.1492,5979.3,2636.4,3351.5,1962.8,0.0000,-7768.7,-7340.2,-1782.4,-2708.5,-3309.4,-17152.,-171.91,-20692.,-6450.5,-4494.3,-2969.5,68.974,2457.1,2240.5,1757.6,346.70,3861.6,1686.6,0.0000,7145.0,4449.7,4252.8,3658.0,0.0000,-404.79,-128.04,-95.612,-45.982,-146.50,-587.69,0.0000,-1087.2,-1615.2,-758.30,-1312.7
584.0000000000,98.698,2052.2,2125.1,1674.6,316.02,3539.5,973.00,1.1498,5974.6,2636.6,3351.5,1963.1,0.0000,-7764.9,-7338.8,-1781.5,-2707.1,-3306.5,-17149.,-171.71,-20689.,-6450.1,-4493.6,-2968.6,68.827,2451.9,2235.8,1750.2,345.89,3844.1,1686.6,0.0000,7134.3,4449.7,4252.8,3658.0,0.0000,-403.84,-127.72,-95.283,-45.885,-145.76,-587.69,0.0000,-1087.0,-1615.0,-758.28,-1312.5
585.0000000000,98.650,2049.8,2123.0,1670.7,315.45,3528.6,972.98,1.1503,5970.7,2636.8,3351.5,1963.3,0.0000,-7760.8,-7337.3,-1780.5,-2705.6,-3303.4,-17146.,-171.50,-20686.,-6449.8,-4492.9,-2967.6,68.652,2445.7,2230.1,1742.5,344.96,3826.1,1686.6,0.0000,7123.4,4449.7,4252.8,3658.0,0.0000,-402.71,-127.35,-94.930,-45.768,-145.00,-587.69,0.0000,-1086.8,-1614.8,-758.27,-1312.2
586.0000000000,98.505,2046.5,2119.9,1665.6,314.69,3520.0,972.97,1.5233,5969.9,2637.0,3351.5,1963.6,0.0000,-7756.4,-7335.6,-1779.3,-2704.1,-3300.1,-17143.,-171.30,-20682.,-6449.4,-4492.2,-2966.6,68.463,2439.0,2223.9,1734.8,343.96,3808.0,1686.6,0.0000,7112.5,4449.7,4252.8,3658.0,0.0000,-401.51,-126.96,-94.567,-45.642,-144.23,-587.69,0.0000,-1086.7,-1614.6,-758.25,-1312.0
587.0000000000,98.327,2042.2,2116.4,1661.3,313.86,3512.8,972.96,1.3805,5967.4,2637.2,3351.6,1963.8,0.0000,-7751.8,-7333.8,-1777.9,-2702.6,-3296.7,-17139.,-171.10,-20679.,-6449.1,-4491.5,-2965.7,68.272,2432.1,2217.7,1727.0,342.95,3790.1,1686.6,0.0000,7101.6,4449.7,4252.8,3658.0,0.0000,-400.28,-126.56,-94.204,-45.515,-143.47,-587.69,0.0000,-1086.5,-1614.5,-758.24,-1311.7
588.0000000000,98.135,2038.5,2112.8,1655.1,312.98,3502.4,972.93,1.5175,5961.8,2637.4,3351.6,1964.1,0.0000,-7747.0,-7331.9,-1776.4,-2701.1,-3293.1,-17136.,-170.90,-20675.,-6448.7,-4490.8,-2964.7,68.073,2425.1,2211.3,1719.2,341.90,3772.0,1686.6,0.0000,7090.6,4449.7,4252.8,3658.0,0.0000,-399.01,-126.14,-93.834,-45.382,-142.70,-587.69,0.0000,-1086.4,-1614.3,-758.22,-1311.5
589.0000000000,97.888,2034.1,2108.1,1649.5,312.18,3489.0,972.94,3.4810,5954.4,2637.6,3351.6,1964.3,0.0000,-7742.2,-7329.9,-1774.9,-2699.6,-3289.4,-17133.,-170.70,-20672.,-6448.3,-4490.1,-2963.7,67.990,2422.1,2208.5,1714.2,341.43,3760.0,1686.6,0.0000,7083.4,4449.7,4252.8,3658.0,0.0000,-398.42,-125.94,-93.620,-45.326,-142.16,-587.69,0.0000,-1086.3,-1614.1,-758.21,-1311.2
590.0000000000,97.681,2031.4,2104.6,1644.0,311.67,3476.7,972.94,3.2082,5946.0,2637.8,3351.4,1964.5,0.0000,-7737.2,-7327.9,-1773.3,-2698.1,-3285.6,-17130.,-170.50,-20668.,-6448.0,-4489.4,-2962.8,68.100,2423.6,2209.5,1711.1,341.52,3751.6,1686.6,97.281,7078.3,4460.9,4252.8,3662.6,0.0000,-398.50,-125.94,-93.530,-45.347,-141.76,-587.69,-4.4556,-1086.2,-1613.9,-758.19,-1311.2
591.0000000000,97.372,2030.3,2102.5,1638.6,311.25,3466.0,972.94,4.0832,5937.6,2638.0,3351.4,1964.8,0.0000,-7732.2,-7326.0,-1771.7,-2696.6,-3281.8,-17127.,-170.31,-20664.,-6447.6,-4488.7,-2961.8,67.824,2416.2,2203.2,1703.4,340.48,3733.7,1686.6,0.0000,7067.4,4449.7,4252.8,3658.0,0.0000,-397.24,-125.53,-93.164,-45.216,-140.99,-587.69,0.0000,-1086.0,-1613.7,-758.18,-1310.8
592.0000000000,97.170,2026.6,2099.1,1633.2,310.59,3453.8,972.94,3.1795,5929.7,2638.2,3351.4,1965.0,0.0000,-7727.1,-7324.0,-1770.1,-2695.1,-3278.0,-17124.,-170.11,-20661.,-6447.2,-4488.0,-2960.8,67.623,2409.0,2196.6,1695.5,339.43,3715.5,1686.6,0.0000,7056.4,4449.7,4252.8,3658.0,0.0000,-395.96,-125.11,-92.791,-45.082,-140.21,-587.69,0.0000,-1085.8,-1613.5,-758.16,-1310.5
593.0000000000,97.024,2021.8,2094.2,1627.4,309.88,3440.5,972.94,3.1817,5921.6,2638.4,3351.4,1965.2,0.0000,-7721.7,-7322.0,-1768.4,-2693.5,-3274.0,-17121.,-169.91,-20657.,-6446.9,-4487.3,-2959.8,67.420,2401.8,2190.0,1687.6,338.36,3697.1,1686.6,0.0000,7045.3,4449.7,4252.8,3658.0,0.0000,-394.66,-124.68,-92.415,-44.946,-139.42,-587.69,0.0000,-1085.7,-1613.3,-758.15,-1310.3
594.0000000000,96.844,2017.1,2089.9,1621.0,309.02,3426.5,972.94,4.1725,5912.7,2638.3,3351.4,1965.5,0.0000,-7716.2,-7319.9,-1766.7,-2692.0,-3269.9,-17118.,-169.72,-20653.,-6446.5,-4486.6,-2958.9,67.306,2397.7,2186.3,1681.1,337.73,3681.7,1686.6,0.0000,7035.9,4449.7,4252.8,3658.0,0.0000,-393.88,-124.41,-92.136,-44.870,-138.74,-587.69,0.0000,-1085.5,-1613.1,-758.14,-1310.1
595.0000000000,96.693,2015.4,2088.2,1614.6,308.74,3412.8,972.94,5.2729,5904.6,2638.5,3351.4,1965.7,0.0000,-7710.9,-7317.9,-1765.0,-2690.4,-3265.8,-17115.,-169.52,-20649.,-6446.1,-4485.9,-2957.9,80.158,2417.4,2209.5,1682.9,341.80,3682.7,1686.6,0.0000,7036.6,4449.7,4257.5,3663.8,0.0000,-395.88,-125.27,-92.360,-45.125,-138.62,-587.69,0.0000,-1085.5,-1613.0,-758.15,-1310.1
596.0000000000,96.809,2020.6,2091.7,1609.5,309.47,3401.6,972.94,5.2733,5899.3,2638.7,3351.4,1965.9,0.0000,-7706.2,-7316.2,-1763.3,-2689.0,-3261.7,-17112.,-169.33,-20644.,-6445.8,-4485.2,-2956.9,123.03,2429.8,2213.0,1680.9,341.49,3671.8,1686.6,0.0000,7029.8,4449.7,4252.8,3658.0,0.0000,-398.47,-125.83,-92.549,-45.418,-138.18,-587.69,0.0000,-1085.4,-1612.8,-758.11,-1309.6
597.0000000000,97.229,2027.4,2097.7,1605.6,310.38,3391.6,972.94,5.2735,5894.2,2638.7,3351.5,1966.1,0.0000,-7702.1,-7314.9,-1761.6,-2687.6,-3257.5,-17108.,-169.13,-20640.,-6445.4,-4484.5,-2955.9,68.193,2429.3,2215.1,1674.4,341.68,3654.2,1686.6,0.0000,7019.0,4449.7,4252.8,3658.0,0.0000,-398.76,-125.92,-92.361,-45.462,-137.42,-587.69,0.0000,-1085.2,-1612.6,-758.09,-1309.4
598.0000000000,97.370,2030.5,2100.5,1603.8,310.91,3380.0,972.94,5.2739,5886.9,2638.9,3351.5,1966.3,0.0000,-7698.2,-7313.7,-1759.9,-2686.2,-3253.4,-17105.,-168.94,-20636.,-6445.0,-4483.8,-2955.0,68.141,2427.5,2213.4,1667.2,341.32,3636.0,1686.6,0.0000,7008.0,4449.7,4252.8,3658.0,0.0000,-398.36,-125.78,-92.087,-45.427,-136.63,-587.69,0.0000,-1085.1,-1612.4,-758.08,-1309.2
599.0000000000,97.482,2030.2,2100.2,1600.8,310.96,3366.6,972.94,5.2741,5878.6,2638.9,3351.5,1966.5,0.0000,-7694.2,-7312.5,-1758.2,-2684.8,-3249.1,-17102.,-168.74,-20632.,-6444.6,-4483.1,-2954.0,68.032,2423.6,2209.9,1659.6,340.69,3617.7,1686.6,0.0000,6996.9,4449.7,4252.8,3658.0,0.0000,-397.63,-125.54,-91.773,-45.355,-135.84,-587.69,0.0000,-1084.9,-1612.2,-758.06,-1309.0
600.0000000000,97.477,2028.5,2098.4,1595.3,310.55,3352.3,972.94,5.2744,5870.9,2639.2,3351.5,1966.8,0.0000,-7690.1,-7311.1,-1756.4,-2683.4,-3244.7,-17099.,-168.55,-20628.,-6444.3,-4482.4,-2953.0,67.894,2418.7,2205.4,1652.0,339.93,3599.5,1686.6,0.0000,6985.8,4449.7,4252.8,3658.0,0.0000,-396.73,-125.24,-91.441,-45.262,-135.04,-587.69,0.0000,-1084.8,-1612.0,-758.05,-1308.7
601.0000000000,97.375,2025.8,2095.5,1589.3,309.94,3337.8,972.94,5.2747,5864.1,2639.5,3351.5,1967.0,0.0000,-7685.7,-7309.5,-1754.5,-2682.0,-3240.2,-17096.,-168.35,-20623.,-6443.9,-4481.7,-2952.0,67.738,2413.1,2200.4,1644.4,339.08,3581.3,1686.6,0.0000,6974.8,4449.7,4252.8,3658.0,0.0000,-395.72,-124.91,-91.099,-45.159,-134.26,-587.69,0.0000,-1084.6,-1611.8,-758.03,-1308.5
602.0000000000,97.234,2021.7,2092.5,1582.7,309.23,3324.5,972.93,5.2750,5857.0,2639.4,3351.6,1967.3,0.0000,-7681.2,-7307.9,-1752.6,-2680.5,-3235.5,-17093.,-168.16,-20619.,-6443.5,-4481.0,-2951.1,67.567,2407.0,2194.8,1636.6,338.16,3563.1,1686.6,0.0000,6963.7,4449.7,4252.8,3658.0,0.0000,-394.63,-124.55,-90.745,-45.045,-133.46,-587.69,0.0000,-1084.5,-1611.7,-758.02,-1308.3
603.0000000000,97.070,2018.0,2089.7,1575.8,308.45,3311.2,972.90,5.8121,5849.5,2639.6,3351.7,1967.5,0.0000,-7676.5,-7306.2,-1750.6,-2679.1,-3230.8,-17090.,-167.97,-20614.,-6443.1,-4480.3,-2950.1,67.389,2400.7,2189.0,1628.8,337.21,3544.9,1686.6,0.0000,6952.7,4449.7,4252.8,3658.0,0.0000,-393.49,-124.18,-90.388,-44.926,-132.67,-587.69,0.0000,-1084.3,-1611.5,-758.00,-1308.1
604.0000000000,96.893,2014.1,2086.1,1569.2,307.64,3296.9,972.90,6.0235,5840.5,2639.8,3351.7,1967.7,0.0000,-7671.7,-7304.3,-1748.5,-2677.6,-3226.1,-17087.,-167.77,-20609.,-6442.7,-4479.6,-2949.1,67.205,2394.2,2183.1,1621.1,336.24,3526.8,1686.6,0.0000,6941.7,4449.7,4252.8,3658.0,0.0000,-392.32,-123.79,-90.028,-44.804,-131.88,-587.69,0.0000,-1084.1,-1611.3,-757.99,-1307.8
605.0000000000,96.708,2009.6,2081.3,1562.7,306.79,3284.4,972.90,5.3004,5831.0,2640.0,3351.6,1967.9,0.0000,-7666.8,-7302.4,-1746.4,-2676.1,-3221.2,-17084.,-167.58,-20605.,-6442.3,-4478.9,-2948.1,67.020,2387.6,2177.1,1613.4,335.25,3508.9,1686.6,0.0000,6930.9,4449.7,4252.8,3658.0,0.0000,-391.13,-123.40,-89.669,-44.680,-131.10,-587.69,0.0000,-1084.0,-1611.1,-757.97,-1307.6
606.0000000000,96.518,2005.0,2076.3,1556.0,305.94,3268.6,972.90,5.3007,5821.3,2640.3,3351.6,1968.2,0.0000,-7661.6,-7300.4,-1744.3,-2674.6,-3216.3,-17081.,-167.38,-20600.,-6441.9,-4478.2,-2947.1,66.833,2380.9,2171.0,1605.7,334.27,3491.0,1686.6,0.0000,6920.1,4449.7,4252.8,3658.0,0.0000,-389.94,-123.00,-89.310,-44.556,-130.31,-587.69,0.0000,-1083.8,-1610.9,-757.96,-1307.4
607.0000000000,96.325,2000.4,2072.1,1549.1,305.12,3253.2,972.90,5.3008,5811.5,2640.7,3351.6,1968.4,0.0000,-7656.2,-7298.3,-1742.1,-2673.0,-3211.3,-17077.,-167.19,-20595.,-6441.6,-4477.5,-2946.2,66.698,2376.1,2166.6,1598.9,333.53,3474.9,1686.6,0.0000,6910.3,4449.7,4252.8,3658.0,0.0000,-389.04,-122.70,-89.008,-44.465,-129.60,-587.69,0.0000,-1083.7,-1610.7,-757.94,-1307.2
608.0000000000,96.158,1996.1,2068.1,1542.2,304.35,3238.1,972.90,5.9943,5802.0,2641.2,3351.6,1968.7,0.0000,-7650.8,-7296.2,-1739.9,-2671.5,-3206.2,-17074.,-167.00,-20590.,-6441.2,-4476.8,-2945.2,66.514,2369.5,2160.6,1591.3,332.55,3457.3,1686.6,0.0000,6899.6,4449.7,4252.8,3658.0,0.0000,-387.86,-122.31,-88.653,-44.343,-128.82,-587.69,0.0000,-1083.5,-1610.5,-757.93,-1307.0
609.0000000000,95.970,1991.2,2063.2,1535.4,303.50,3225.9,972.90,7.1720,5792.4,2641.4,3351.6,1968.9,0.0000,-7645.2,-7294.0,-1737.7,-2670.0,-3201.1,-17071.,-166.81,-20585.,-6440.8,-4476.1,-2944.2,66.295,2361.7,2153.5,1583.0,331.41,3438.2,1686.6,0.0000,6888.1,4449.7,4252.8,3658.0,0.0000,-386.47,-121.85,-88.257,-44.196,-127.99,-587.69,0.0000,-1083.4,-1610.4,-757.91,-1306.7
610.0000000000,95.767,1985.7,2057.8,1528.4,302.59,3211.1,972.90,5.3596,5782.9,2641.6,3351.7,1969.1,0.0000,-7639.4,-7291.7,-1735.4,-2668.4,-3196.0,-17068.,-166.61,-20581.,-6440.4,-4475.4,-2943.2,66.074,2353.9,2146.3,1574.8,330.25,3419.2,1686.6,0.0000,6876.6,4449.7,4252.8,3658.0,0.0000,-385.07,-121.39,-87.861,-44.050,-127.16,-587.69,0.0000,-1083.2,-1610.2,-757.90,-1306.5
611.0000000000,95.557,1979.9,2052.0,1521.1,301.63,3195.1,972.90,5.3598,5773.3,2641.7,3351.7,1969.3,0.0000,-7633.5,-7289.4,-1733.1,-2666.9,-3190.7,-17065.,-166.42,-20576.,-6440.0,-4474.7,-2942.2,65.863,2346.3,2139.5,1566.7,329.14,3400.7,1686.6,0.0000,6865.4,4449.7,4252.8,3658.0,0.0000,-383.72,-120.94,-87.477,-43.909,-126.35,-587.69,0.0000,-1083.0,-1610.0,-757.88,-1306.3
612.0000000000,95.252,1974.2,2046.1,1513.7,300.67,3179.2,972.86,5.3600,5763.8,2641.9,3351.8,1969.5,0.0000,-7627.4,-7287.0,-1730.7,-2665.3,-3185.4,-17062.,-166.23,-20571.,-6439.7,-4473.9,-2941.3,65.675,2339.6,2133.4,1558.9,328.15,3382.7,1686.6,0.0000,6854.4,4449.7,4252.8,3658.0,0.0000,-382.51,-120.54,-87.115,-43.784,-125.56,-587.69,0.0000,-1082.9,-1609.8,-757.87,-1306.1
613.0000000000,94.847,1969.3,2041.0,1506.6,299.86,3163.9,972.86,5.3602,5754.3,2642.1,3351.7,1969.7,0.0000,-7621.3,-7284.5,-1728.4,-2663.8,-3180.0,-17059.,-166.04,-20565.,-6439.3,-4473.2,-2940.3,65.617,2337.6,2132.2,1559.0,328.94,3382.9,1686.6,6.9868,6855.3,4452.9,4255.7,3661.8,0.0000,-382.05,-120.39,-87.066,-43.751,-125.43,-587.69,-0.32000,-1082.9,-1609.6,-757.87,-1306.0
614.0000000000,94.712,1966.0,2037.2,1500.6,299.33,3150.5,972.86,5.3604,5745.3,2642.3,3351.8,1969.9,0.0000,-7615.1,-7282.1,-1726.0,-2662.2,-3174.7,-17056.,-165.85,-20560.,-6438.9,-4472.5,-2939.3,65.553,2335.3,2129.4,1552.1,327.47,3366.2,1686.6,0.0000,6844.4,4449.7,4252.8,3658.0,0.0000,-381.56,-120.20,-86.817,-43.702,-124.72,-587.69,0.0000,-1082.7,-1609.4,-757.84,-1305.6
615.0000000000,94.594,1962.8,2033.6,1495.3,298.82,3137.6,972.86,5.3607,5736.8,2642.5,3351.8,1970.2,0.0000,-7609.1,-7279.8,-1723.7,-2660.7,-3169.3,-17052.,-165.66,-20555.,-6438.5,-4471.8,-2938.3,65.365,2328.6,2123.3,1544.6,326.48,3348.9,1686.6,0.0000,6833.9,4449.7,4252.8,3658.0,0.0000,-380.34,-119.79,-86.463,-43.576,-123.95,-587.69,0.0000,-1082.6,-1609.3,-757.82,-1305.4
616.0000000000,94.442,1959.9,2030.3,1489.9,298.40,3124.0,972.86,5.3609,5728.0,2642.7,3351.8,1970.4,0.0000,-7603.0,-7277.4,-1721.4,-2659.1,-3164.0,-17049.,-165.48,-20550.,-6438.1,-4471.1,-2937.4,68.022,2333.2,2128.9,1542.1,327.02,3341.0,1686.6,0.0000,6829.1,4449.7,4252.8,3658.0,0.0000,-380.97,-120.00,-86.444,-43.662,-123.54,-587.69,0.0000,-1082.5,-1609.1,-757.81,-1305.2
617.0000000000,94.453,1958.6,2028.2,1484.8,298.26,3110.6,972.82,5.3611,5719.2,2642.9,3351.8,1970.7,0.0000,-7597.1,-7275.2,-1719.1,-2657.6,-3158.7,-17046.,-165.29,-20545.,-6437.8,-4470.4,-2936.4,65.327,2327.3,2122.1,1534.6,326.14,3323.5,1686.6,0.0000,6818.5,4449.7,4252.8,3658.0,0.0000,-379.89,-119.61,-86.104,-43.552,-122.76,-587.69,0.0000,-1082.3,-1608.9,-757.79,-1305.0
618.0000000000,94.329,1955.5,2025.4,1479.5,297.60,3097.0,972.82,5.3614,5710.6,2643.1,3351.8,1970.9,0.0000,-7591.2,-7272.9,-1716.8,-2656.1,-3153.2,-17043.,-165.10,-20540.,-6437.4,-4469.7,-2935.4,65.147,2320.8,2116.2,1527.0,325.18,3305.7,1686.6,0.0000,6807.7,4449.7,4252.8,3658.0,0.0000,-378.73,-119.22,-85.751,-43.432,-121.98,-587.69,0.0000,-1082.2,-1608.7,-757.78,-1304.8
619.0000000000,94.196,1951.2,2021.3,1473.8,296.98,3082.7,972.82,4.4992,5702.1,2643.1,3351.8,1971.1,0.0000,-7585.2,-7270.6,-1714.5,-2654.5,-3147.8,-17040.,-164.91,-20535.,-6437.0,-4469.0,-2934.4,64.959,2314.1,2110.1,1519.4,324.19,3287.9,1686.6,0.0000,6797.0,4449.7,4252.8,3658.0,0.0000,-377.51,-118.82,-85.392,-43.306,-121.19,-587.69,0.0000,-1082.0,-1608.5,-757.76,-1304.6
620.0000000000,94.053,1946.4,2017.1,1467.4,296.16,3069.1,972.82,5.4252,5694.4,2643.3,3351.8,1971.3,0.0000,-7579.0,-7268.2,-1712.1,-2653.0,-3142.2,-17037.,-164.72,-20529.,-6436.6,-4468.2,-2933.4,64.791,2308.1,2104.6,1512.1,323.29,3271.0,1686.6,0.0000,6786.7,4449.7,4252.8,3658.0,0.0000,-376.42,-118.45,-85.057,-43.194,-120.44,-587.69,0.0000,-1081.8,-1608.4,-757.75,-1304.3
621.0000000000,93.873,1942.1,2012.7,1460.7,295.40,3055.7,972.82,5.4254,5686.4,2643.6,3351.8,1971.5,0.0000,-7572.8,-7265.7,-1709.7,-2651.4,-3136.6,-17034.,-164.53,-20524.,-6436.2,-4467.5,-2932.5,64.687,2304.4,2101.3,1506.4,322.71,3257.4,1686.6,0.0000,6778.4,4449.7,4252.8,3658.0,0.0000,-375.69,-118.20,-84.808,-43.125,-119.81,-587.69,0.0000,-1081.7,-1608.2,-757.73,-1304.1
622.0000000000,93.726,1938.8,2009.2,1454.6,294.76,3042.1,972.82,5.4256,5678.0,2643.8,3351.9,1971.7,0.0000,-7566.7,-7263.3,-1707.3,-2649.9,-3131.0,-17030.,-164.35,-20519.,-6435.8,-4466.8,-2931.5,64.634,2302.5,2099.5,1501.8,322.39,3246.0,1686.6,0.0000,6771.5,4449.7,4252.8,3658.0,0.0000,-375.26,-118.04,-84.623,-43.089,-119.27,-587.69,0.0000,-1081.6,-1608.0,-757.72,-1303.9
623.0000000000,93.615,1935.7,2006.3,1448.8,294.23,3029.1,972.82,4.1148,5670.0,2644.2,3351.9,1971.9,0.0000,-7560.6,-7260.9,-1704.8,-2648.3,-3125.3,-17027.,-164.16,-20514.,-6435.4,-4466.1,-2930.5,64.486,2297.3,2094.8,1495.3,321.60,3230.7,1686.6,0.0000,6762.2,4449.7,4252.8,3658.0,0.0000,-374.29,-117.71,-84.324,-42.991,-118.58,-587.69,0.0000,-1081.5,-1607.8,-757.70,-1303.7
624.0000000000,93.476,1932.2,2002.7,1443.1,293.62,3016.1,972.82,3.4658,5661.6,2644.4,3351.9,1972.1,0.0000,-7554.4,-7258.5,-1702.4,-2646.8,-3119.7,-17024.,-163.97,-20508.,-6435.0,-4465.4,-2929.5,64.324,2291.5,2089.5,1488.4,320.74,3214.5,1686.6,0.0000,6752.5,4449.7,4252.8,3658.0,0.0000,-373.22,-117.35,-84.003,-42.882,-117.85,-587.69,0.0000,-1081.3,-1607.6,-757.69,-1303.5
625.0000000000,93.335,1928.4,1998.5,1437.2,293.02,3002.3,972.82,3.4661,5652.7,2644.3,3351.9,1972.3,0.0000,-7548.2,-7256.1,-1699.9,-2645.2,-3114.0,-17021.,-163.79,-20503.,-6434.6,-4464.6,-2928.6,64.205,2287.3,2085.6,1482.2,320.09,3199.9,1686.6,0.0000,6743.6,4449.7,4252.8,3658.0,0.0000,-372.41,-117.08,-83.732,-42.803,-117.18,-587.69,0.0000,-1081.2,-1607.5,-757.67,-1303.3
626.0000000000,93.207,1924.5,1994.3,1431.3,292.36,2988.4,972.82,3.4664,5643.9,2644.4,3351.9,1972.5,0.0000,-7541.9,-7253.6,-1697.5,-2643.7,-3108.2,-17018.,-163.60,-20497.,-6434.2,-4463.9,-2927.6,64.037,2281.3,2080.1,1475.2,319.20,3183.7,1686.6,0.0000,6733.7,4449.7,4252.8,3658.0,0.0000,-371.32,-116.71,-83.406,-42.691,-116.46,-587.69,0.0000,-1081.0,-1607.3,-757.65,-1303.0
627.0000000000,93.044,1921.3,1990.8,1425.3,291.79,2974.8,972.82,3.4668,5635.4,2644.4,3352.0,1972.7,0.0000,-7535.7,-7251.2,-1695.0,-2642.1,-3102.5,-17015.,-163.42,-20492.,-6433.8,-4463.2,-2926.6,64.096,2283.4,2082.1,1474.1,319.45,3180.7,1686.6,10.400,6733.5,4454.1,4256.9,3662.9,0.0000,-371.54,-116.76,-83.389,-42.731,-116.18,-587.69,-0.47634,-1081.0,-1607.1,-757.66,-1303.0
628.0000000000,92.996,1919.3,1988.5,1420.0,291.51,2962.4,972.82,3.4671,5627.3,2644.6,3352.0,1972.9,0.0000,-7529.5,-7248.8,-1692.6,-2640.6,-3096.7,-17011.,-163.23,-20487.,-6433.4,-4462.5,-2925.6,63.955,2278.4,2077.5,1468.1,318.70,3166.1,1686.6,0.0000,6723.1,4449.8,4253.0,3659.5,0.0000,-370.60,-116.44,-83.120,-42.637,-115.56,-587.69,0.0000,-1080.8,-1606.9,-757.62,-1302.7
629.0000000000,92.875,1917.1,1986.3,1415.3,291.09,2954.7,972.79,3.4674,5619.6,2644.8,3352.0,1973.1,0.0000,-7523.4,-7246.5,-1690.2,-2639.0,-3091.0,-17008.,-163.05,-20481.,-6433.0,-4461.7,-2924.7,63.978,2279.6,2078.3,1471.6,321.12,3173.3,1686.6,20.239,6726.0,4453.0,4252.9,3658.6,0.0000,-370.62,-116.43,-83.194,-42.666,-115.62,-587.69,-0.92694,-1080.8,-1606.7,-757.61,-1302.4
630.0000000000,92.841,1916.5,1985.2,1411.4,291.13,2945.7,972.78,3.4677,5612.7,2644.9,3352.0,1973.3,0.0000,-7517.5,-7244.3,-1687.8,-2637.5,-3085.3,-17005.,-162.87,-20476.,-6432.6,-4461.0,-2923.7,64.076,2284.3,2082.3,1467.5,319.80,3163.0,1686.6,0.0000,6721.2,4449.7,4252.8,3658.4,0.0000,-371.07,-116.56,-83.160,-42.721,-115.21,-587.69,0.0000,-1080.7,-1606.6,-757.59,-1302.2
631.0000000000,92.874,1916.5,1984.8,1408.6,291.12,2936.8,972.78,3.4680,5605.7,2645.1,3352.1,1973.6,0.0000,-7511.8,-7242.2,-1685.5,-2636.0,-3079.8,-17002.,-162.69,-20471.,-6432.2,-4460.3,-2922.7,63.968,2278.8,2077.9,1461.2,318.64,3148.1,1686.6,0.0000,6712.1,4449.7,4252.8,3658.3,0.0000,-370.33,-116.29,-82.891,-42.645,-114.53,-587.69,0.0000,-1080.6,-1606.4,-757.58,-1302.0
632.0000000000,92.801,1914.8,1982.9,1405.1,290.82,2926.7,972.78,3.4684,5599.1,2645.3,3352.1,1973.8,0.0000,-7506.1,-7240.1,-1683.2,-2634.6,-3074.2,-16999.,-162.50,-20466.,-6431.8,-4459.6,-2921.7,63.845,2274.4,2073.9,1454.9,317.97,3133.1,1686.6,0.0000,6703.0,4449.7,4252.8,3658.1,0.0000,-369.50,-116.01,-82.612,-42.563,-113.86,-587.69,0.0000,-1080.5,-1606.2,-757.56,-1301.8
633.0000000000,92.733,1912.1,1980.1,1401.3,290.46,2915.2,972.78,3.2001,5591.9,2645.5,3352.1,1974.0,0.0000,-7500.3,-7238.0,-1680.9,-2633.1,-3068.6,-16996.,-162.32,-20460.,-6431.4,-4458.8,-2920.7,63.735,2270.5,2070.3,1449.0,317.36,3119.0,1686.6,0.0000,6694.5,4449.7,4252.8,3658.0,0.0000,-368.75,-115.76,-82.353,-42.490,-113.21,-587.69,0.0000,-1080.3,-1606.0,-757.54,-1301.5
634.0000000000,92.649,1909.2,1977.4,1396.4,289.90,2903.6,972.82,1.4251,5585.4,2645.6,3352.1,1974.2,0.0000,-7494.5,-7235.9,-1678.6,-2631.6,-3062.9,-16993.,-162.14,-20455.,-6431.0,-4458.1,-2919.8,63.610,2266.1,2066.3,1443.1,316.69,3104.9,1686.6,0.0000,6685.9,4449.7,4252.8,3658.0,0.0000,-367.92,-115.48,-82.086,-42.407,-112.57,-587.69,0.0000,-1080.2,-1605.8,-757.53,-1301.3
635.0000000000,92.536,1912.6,1980.5,1392.0,290.46,2894.0,972.86,1.4256,5579.2,2645.7,3352.0,1974.4,0.0000,-7489.2,-7234.0,-1676.4,-2630.1,-3057.2,-16989.,-161.96,-20450.,-6430.6,-4457.4,-2918.8,69.670,2326.9,2118.5,1469.1,332.60,3150.7,1686.6,161.49,6716.4,4463.5,4263.4,3672.5,0.0000,-375.37,-118.01,-83.448,-43.335,-113.90,-587.69,-7.3966,-1080.5,-1605.7,-757.57,-1301.8
636.0000000000,93.157,1928.6,1993.5,1390.5,293.01,2890.3,972.83,1.4262,5575.6,2645.9,3352.0,1974.6,0.0000,-7485.2,-7232.9,-1674.3,-2628.8,-3051.7,-16986.,-161.78,-20445.,-6430.1,-4456.6,-2917.8,65.379,2343.8,2140.8,1471.5,336.44,3151.3,1686.6,36.334,6716.7,4467.8,4266.8,3682.7,0.0000,-377.98,-118.97,-83.763,-43.657,-113.79,-587.69,-1.6641,-1080.5,-1605.5,-757.57,-1302.0
637.0000000000,93.538,1941.7,2006.8,1392.2,294.64,2889.6,972.81,1.5026,5572.5,2645.9,3352.0,1974.8,0.0000,-7482.2,-7232.3,-1672.4,-2627.6,-3046.4,-16983.,-161.60,-20440.,-6429.7,-4455.9,-2916.9,65.591,2336.7,2130.6,1462.4,326.16,3132.9,1686.6,0.0000,6703.1,4458.7,4258.7,3670.4,0.0000,-379.10,-118.96,-83.763,-43.728,-113.23,-587.69,0.0000,-1080.3,-1605.3,-757.51,-1301.3
638.0000000000,93.862,1949.3,2014.2,1393.0,296.42,2886.4,972.81,1.5048,5568.8,2645.9,3352.0,1975.0,0.0000,-7479.4,-7231.7,-1670.5,-2626.4,-3041.3,-16980.,-161.42,-20435.,-6429.3,-4455.2,-2915.9,65.602,2337.0,2131.0,1457.3,326.09,3119.5,1686.6,0.0000,6694.6,4453.9,4255.5,3663.9,0.0000,-379.09,-118.95,-83.595,-43.735,-112.62,-587.69,0.0000,-1080.1,-1605.1,-757.48,-1300.8
639.0000000000,93.932,1952.2,2017.5,1392.9,296.93,2879.6,972.76,1.5054,5563.5,2646.0,3352.1,1975.2,0.0000,-7476.7,-7231.1,-1668.6,-2625.1,-3036.0,-16977.,-161.24,-20430.,-6428.9,-4454.4,-2914.9,65.529,2334.4,2128.6,1451.4,325.64,3104.8,1686.6,0.0000,6685.6,4451.0,4253.7,3659.8,0.0000,-378.59,-118.79,-83.355,-43.686,-111.97,-587.69,0.0000,-1080.0,-1605.0,-757.45,-1300.4
640.0000000000,93.721,1952.5,2018.3,1390.5,296.84,2870.7,972.73,1.5060,5558.3,2646.0,3352.1,1975.5,0.0000,-7473.7,-7230.3,-1666.6,-2623.9,-3030.7,-16974.,-161.06,-20425.,-6428.5,-4453.7,-2913.9,65.410,2330.2,2124.8,1445.0,324.98,3089.7,1686.6,0.0000,6676.3,4450.0,4253.0,3658.4,0.0000,-377.83,-118.54,-83.077,-43.607,-111.29,-587.69,0.0000,-1079.9,-1604.8,-757.43,-1300.1
641.0000000000,93.674,1951.5,2017.1,1387.4,296.42,2860.0,972.73,1.5065,5552.8,2646.2,3352.1,1975.7,0.0000,-7470.4,-7229.4,-1664.7,-2622.6,-3025.2,-16970.,-160.88,-20420.,-6428.1,-4453.0,-2913.0,65.297,2326.2,2121.1,1439.1,324.36,3075.5,1686.6,0.0000,6667.7,4449.7,4252.8,3658.0,0.0000,-377.11,-118.31,-82.815,-43.531,-110.65,-587.69,0.0000,-1079.7,-1604.6,-757.42,-1299.9
642.0000000000,93.577,1949.5,2016.1,1382.6,295.91,2850.6,972.70,1.5071,5550.1,2646.4,3352.1,1975.9,0.0000,-7466.9,-7228.3,-1662.6,-2621.3,-3019.6,-16967.,-160.70,-20415.,-6427.7,-4452.2,-2912.0,65.185,2322.2,2117.5,1433.3,323.75,3061.9,1686.6,0.0000,6659.4,4449.7,4252.8,3658.0,0.0000,-376.39,-118.07,-82.561,-43.457,-110.03,-587.69,0.0000,-1079.6,-1604.5,-757.40,-1299.7
643.0000000000,93.461,1947.8,2014.9,1377.2,295.36,2843.9,972.68,1.5076,5547.6,2646.5,3352.1,1976.1,0.0000,-7463.4,-7227.2,-1660.4,-2619.9,-3014.0,-16964.,-160.52,-20410.,-6427.2,-4451.5,-2911.0,65.066,2318.0,2113.6,1427.6,323.11,3048.2,1686.6,0.0000,6651.2,4449.7,4252.8,3658.0,0.0000,-375.63,-117.82,-82.303,-43.378,-109.41,-587.69,0.0000,-1079.5,-1604.3,-757.39,-1299.5
644.0000000000,93.336,1945.6,2012.7,1372.3,294.78,2840.1,972.65,1.5082,5543.7,2646.7,3352.1,1976.3,0.0000,-7459.7,-7225.9,-1658.2,-2618.6,-3008.4,-16961.,-160.34,-20405.,-6426.8,-4450.7,-2910.0,64.924,2312.9,2109.0,1421.5,322.35,3034.0,1686.6,0.0000,6642.6,4449.7,4252.8,3658.0,0.0000,-374.73,-117.53,-82.022,-43.283,-108.77,-587.69,0.0000,-1079.3,-1604.1,-757.37,-1299.3
645.0000000000,93.198,1942.4,2009.1,1367.9,294.15,2830.7,972.65,1.5088,5538.2,2646.9,3352.1,1976.5,0.0000,-7455.8,-7224.5,-1655.9,-2617.2,-3002.7,-16958.,-160.16,-20400.,-6426.4,-4450.0,-2909.1,64.774,2307.5,2104.1,1415.4,321.55,3019.8,1686.6,0.0000,6633.9,4449.7,4252.8,3658.0,0.0000,-373.79,-117.22,-81.734,-43.182,-108.13,-587.69,0.0000,-1079.2,-1603.9,-757.35,-1299.1
646.0000000000,93.052,1939.5,2005.2,1363.0,293.49,2819.3,972.65,1.5123,5531.5,2647.1,3352.1,1976.8,0.0000,-7451.7,-7223.1,-1653.6,-2615.8,-2997.0,-16955.,-159.98,-20396.,-6426.0,-4449.3,-2908.1,64.621,2302.1,2099.1,1409.2,320.75,3005.6,1686.6,0.0000,6625.3,4449.7,4252.8,3658.0,0.0000,-372.83,-116.90,-81.446,-43.080,-107.48,-587.69,0.0000,-1079.1,-1603.8,-757.34,-1298.9
647.0000000000,92.899,1936.3,2001.6,1357.7,292.79,2806.9,972.64,1.5225,5524.2,2647.3,3352.1,1977.0,0.0000,-7447.3,-7221.6,-1651.2,-2614.5,-2991.2,-16951.,-159.80,-20391.,-6425.5,-4448.5,-2907.1,64.467,2296.6,2094.1,1403.1,319.94,2991.5,1686.6,0.0000,6616.8,4449.7,4252.8,3658.0,0.0000,-371.86,-116.59,-81.158,-42.978,-106.85,-587.69,0.0000,-1078.9,-1603.6,-757.32,-1298.7
648.0000000000,92.740,1932.4,1997.7,1352.2,292.09,2794.2,972.64,1.5231,5516.5,2647.5,3352.1,1977.2,0.0000,-7442.7,-7220.0,-1648.9,-2613.1,-2985.5,-16948.,-159.62,-20386.,-6425.1,-4447.8,-2906.1,64.312,2291.1,2089.1,1397.1,319.12,2977.5,1686.6,0.0000,6608.3,4449.7,4252.8,3658.0,0.0000,-370.88,-116.26,-80.871,-42.874,-106.21,-587.69,0.0000,-1078.8,-1603.4,-757.30,-1298.5
649.0000000000,92.583,1930.8,1995.8,1346.8,291.76,2783.1,972.64,1.5236,5509.2,2647.9,3352.1,1977.4,0.0000,-7438.2,-7218.4,-1646.5,-2611.7,-2979.7,-16945.,-159.45,-20382.,-6424.7,-4447.0,-2905.2,69.752,2315.2,2114.3,1406.0,330.51,2987.6,1686.6,263.01,6621.1,4470.5,4263.0,3676.9,0.0000,-372.72,-117.13,-81.166,-43.156,-106.33,-587.69,-12.046,-1078.9,-1603.2,-757.34,-1299.1
650.0000000000,92.675,1933.1,1997.8,1342.4,292.08,2773.9,972.67,1.5242,5502.8,2648.2,3352.1,1977.6,0.0000,-7434.1,-7217.1,-1644.2,-2610.4,-2974.0,-16942.,-159.27,-20377.,-6424.3,-4446.3,-2904.2,64.633,2302.5,2099.5,1396.4,320.58,2972.1,1686.6,0.0000,6605.0,4449.7,4252.8,3658.0,0.0000,-372.57,-116.77,-81.012,-43.088,-105.77,-587.69,0.0000,-1078.7,-1603.1,-757.27,-1298.1
651.0000000000,92.656,1933.9,1998.8,1339.5,292.02,2765.6,972.69,1.5248,5496.4,2648.4,3352.1,1977.8,0.0000,-7430.1,-7215.8,-1641.9,-2609.0,-2968.4,-16939.,-159.10,-20373.,-6423.9,-4445.5,-2903.2,64.571,2300.3,2097.5,1391.5,320.22,2960.2,1686.6,0.0000,6597.7,4449.7,4252.8,3658.0,0.0000,-372.13,-116.62,-80.814,-43.047,-105.21,-587.69,0.0000,-1078.6,-1602.9,-757.25,-1297.9
652.0000000000,92.415,1933.2,1997.8,1335.9,292.07,2756.3,972.67,1.5398,5489.8,2648.6,3352.2,1978.0,0.0000,-7426.1,-7214.5,-1639.7,-2607.7,-2962.8,-16936.,-158.92,-20369.,-6423.4,-4444.8,-2902.3,64.511,2298.2,2095.5,1387.0,319.86,2948.9,1686.6,0.0000,6590.9,4449.7,4252.8,3658.0,0.0000,-371.70,-116.47,-80.626,-43.007,-104.68,-587.69,0.0000,-1078.4,-1602.7,-757.24,-1297.7
653.0000000000,92.363,1931.6,1996.2,1332.3,291.82,2746.1,972.67,1.5409,5483.3,2648.7,3352.2,1978.2,0.0000,-7422.0,-7213.2,-1637.4,-2606.4,-2957.2,-16933.,-158.75,-20366.,-6423.0,-4444.0,-2901.3,64.435,2295.4,2093.1,1382.2,319.43,2937.5,1686.6,0.0000,6584.0,4449.7,4252.8,3658.0,0.0000,-371.19,-116.30,-80.425,-42.956,-104.14,-587.69,0.0000,-1078.3,-1602.5,-757.22,-1297.5
654.0000000000,92.294,1929.8,1994.4,1328.3,291.45,2735.6,972.66,1.5415,5477.1,2648.9,3352.2,1978.3,0.0000,-7417.9,-7211.8,-1635.1,-2605.0,-2951.5,-16929.,-158.58,-20362.,-6422.6,-4443.3,-2900.3,64.345,2292.3,2090.2,1377.4,318.93,2925.9,1686.6,0.0000,6577.0,4449.7,4252.8,3658.0,0.0000,-370.59,-116.10,-80.213,-42.897,-103.59,-587.69,0.0000,-1078.2,-1602.4,-757.21,-1297.3
655.0000000000,92.207,1927.5,1991.5,1324.2,291.04,2725.0,972.63,1.5420,5470.7,2649.1,3352.2,1978.5,0.0000,-7413.7,-7210.4,-1632.8,-2603.7,-2945.9,-16926.,-158.40,-20359.,-6422.2,-4442.5,-2899.4,64.241,2288.5,2086.8,1372.4,318.37,2914.1,1686.6,0.0000,6569.8,4449.7,4252.8,3658.0,0.0000,-369.91,-115.87,-79.988,-42.827,-103.04,-587.69,0.0000,-1078.1,-1602.2,-757.19,-1297.1
656.0000000000,92.109,1925.0,1988.7,1319.7,290.57,2715.9,972.63,1.5425,5465.2,2649.3,3352.2,1978.7,0.0000,-7409.4,-7208.8,-1630.5,-2602.3,-2940.2,-16923.,-158.23,-20356.,-6421.8,-4441.8,-2898.4,64.128,2284.5,2083.1,1367.3,317.77,2902.1,1686.6,0.0000,6562.5,4449.7,4252.8,3658.0,0.0000,-369.18,-115.63,-79.755,-42.752,-102.48,-587.69,0.0000,-1078.0,-1602.0,-757.17,-1296.9
657.0000000000,92.108,1922.2,1986.0,1315.2,290.06,2709.0,972.63,1.5431,5460.0,2649.4,3352.3,1978.9,0.0000,-7405.0,-7207.3,-1628.2,-2601.0,-2934.5,-16920.,-158.06,-20353.,-6421.4,-4441.0,-2897.5,64.009,2280.3,2079.2,1362.1,317.13,2890.0,1686.6,0.0000,6555.2,4449.7,4252.8,3658.0,0.0000,-368.41,-115.37,-79.517,-42.672,-101.91,-587.69,0.0000,-1077.8,-1601.9,-757.16,-1296.7
658.0000000000,92.067,1919.3,1983.2,1310.6,289.53,2700.1,972.59,1.5436,5454.3,2649.6,3352.3,1979.0,0.0000,-7400.5,-7205.6,-1625.8,-2599.6,-2928.7,-16917.,-157.88,-20350.,-6420.9,-4440.3,-2896.5,63.892,2276.1,2075.4,1357.0,316.51,2878.2,1686.6,0.0000,6548.0,4449.7,4252.8,3658.0,0.0000,-367.65,-115.12,-79.283,-42.595,-101.36,-587.69,0.0000,-1077.7,-1601.7,-757.14,-1296.5
659.0000000000,91.945,1916.3,1980.9,1306.1,289.02,2690.1,972.59,1.5875,5448.6,2649.8,3352.3,1979.2,0.0000,-7396.0,-7203.9,-1623.5,-2598.2,-2923.0,-16914.,-157.71,-20347.,-6420.5,-4439.5,-2895.5,63.820,2273.6,2073.1,1353.1,316.11,2868.8,1686.6,0.0000,6542.3,4449.7,4252.8,3658.0,0.0000,-367.15,-114.94,-79.112,-42.547,-100.89,-587.69,0.0000,-1077.6,-1601.5,-757.12,-1296.3
660.0000000000,91.845,1914.3,1979.1,1301.6,288.61,2680.0,972.60,1.6225,5442.9,2650.1,3352.3,1979.5,0.0000,-7391.4,-7202.2,-1621.1,-2596.8,-2917.2,-16911.,-157.55,-20344.,-6420.1,-4438.8,-2894.6,63.773,2271.9,2071.6,1349.7,315.84,2860.6,1686.6,0.0000,6537.3,4449.7,4252.8,3658.0,0.0000,-366.80,-114.82,-78.973,-42.515,-100.47,-587.69,0.0000,-1077.5,-1601.3,-757.11,-1296.1
661.0000000000,92.046,1913.8,1978.3,1297.6,288.46,2671.0,972.60,1.6230,5436.7,2650.2,3352.3,1979.6,0.0000,-7387.0,-7200.6,-1618.8,-2595.5,-2911.4,-16907.,-157.38,-20341.,-6419.7,-4438.0,-2893.6,64.870,2281.2,2079.0,1351.7,317.04,2860.8,1686.6,23.698,6539.2,4454.2,4255.2,3662.2,0.0000,-367.82,-115.15,-79.088,-42.644,-100.31,-587.69,-1.0854,-1077.4,-1601.2,-757.10,-1296.1
662.0000000000,92.181,1914.8,1978.6,1294.2,288.60,2662.5,972.60,1.6236,5431.0,2650.4,3352.3,1979.8,0.0000,-7382.8,-7199.1,-1616.5,-2594.2,-2905.7,-16904.,-157.21,-20338.,-6419.3,-4437.3,-2892.6,63.882,2275.8,2075.1,1345.8,316.27,2849.0,1686.6,0.0000,6530.3,4449.7,4252.8,3658.0,0.0000,-367.26,-114.93,-78.893,-42.588,-99.792,-587.69,0.0000,-1077.3,-1601.0,-757.07,-1295.7
663.0000000000,92.137,1914.0,1978.5,1291.3,288.39,2654.4,972.56,1.6255,5425.1,2650.5,3352.3,1980.0,0.0000,-7378.6,-7197.6,-1614.2,-2592.8,-2900.0,-16901.,-157.05,-20335.,-6418.9,-4436.5,-2891.7,63.787,2272.4,2072.0,1341.2,315.75,2838.1,1686.6,0.0000,6523.7,4449.7,4252.8,3658.0,0.0000,-366.63,-114.72,-78.686,-42.525,-99.270,-587.69,0.0000,-1077.1,-1600.8,-757.05,-1295.5
664.0000000000,92.090,1912.0,1977.0,1287.9,288.20,2645.9,972.56,1.6362,5419.4,2650.5,3352.3,1980.2,0.0000,-7374.4,-7196.0,-1611.9,-2591.5,-2894.4,-16898.,-156.88,-20332.,-6418.4,-4435.8,-2890.7,63.687,2268.8,2068.8,1336.5,315.21,2827.1,1686.6,0.0000,6517.0,4449.7,4252.8,3658.0,0.0000,-365.98,-114.50,-78.475,-42.458,-98.747,-587.69,0.0000,-1077.0,-1600.7,-757.04,-1295.3
665.0000000000,92.066,1909.6,1974.7,1284.3,287.76,2636.8,972.54,1.6367,5413.5,2650.7,3352.4,1980.4,0.0000,-7370.1,-7194.4,-1609.6,-2590.1,-2888.7,-16895.,-156.71,-20329.,-6418.0,-4435.0,-2889.7,63.584,2265.1,2065.4,1331.8,314.66,2816.2,1686.6,0.0000,6510.4,4449.7,4252.8,3658.0,0.0000,-365.30,-114.27,-78.262,-42.389,-98.224,-587.69,0.0000,-1076.8,-1600.5,-757.02,-1295.1
666.0000000000,92.123,1907.1,1972.1,1280.3,287.29,2627.4,972.50,1.6373,5407.5,2650.9,3352.4,1980.6,0.0000,-7365.7,-7192.8,-1607.2,-2588.8,-2883.0,-16892.,-156.55,-20326.,-6417.6,-4434.3,-2888.8,63.477,2261.4,2062.0,1327.2,314.09,2805.3,1686.6,0.0000,6503.8,4449.7,4252.8,3658.0,0.0000,-364.61,-114.04,-78.048,-42.318,-97.704,-587.69,0.0000,-1076.7,-1600.3,-757.00,-1294.9
667.0000000000,92.012,1904.2,1969.2,1276.2,286.80,2618.1,972.47,1.6378,5401.8,2651.0,3352.4,1980.8,0.0000,-7361.2,-7191.1,-1604.9,-2587.4,-2877.3,-16889.,-156.38,-20323.,-6417.2,-4433.5,-2887.8,63.373,2257.6,2058.6,1322.6,313.54,2794.5,1686.6,0.0000,6497.3,4449.7,4252.8,3658.0,0.0000,-363.92,-113.81,-77.838,-42.249,-97.190,-587.69,0.0000,-1076.6,-1600.2,-756.99,-1294.7
668.0000000000,91.901,1901.3,1966.4,1271.9,286.31,2608.7,972.47,1.6383,5396.6,2651.2,3352.4,1981.0,0.0000,-7356.7,-7189.4,-1602.6,-2586.1,-2871.5,-16885.,-156.22,-20320.,-6416.8,-4432.8,-2886.8,63.269,2253.9,2055.2,1318.0,312.98,2783.9,1686.6,0.0000,6490.8,4449.7,4252.8,3658.0,0.0000,-363.24,-113.58,-77.628,-42.180,-96.679,-587.69,0.0000,-1076.4,-1600.0,-756.97,-1294.5
669.0000000000,91.789,1898.5,1963.5,1267.5,285.82,2599.7,972.44,1.7151,5391.6,2651.3,3352.4,1981.2,0.0000,-7352.0,-7187.6,-1600.2,-2584.7,-2865.7,-16882.,-156.05,-20318.,-6416.3,-4432.0,-2885.9,63.164,2250.2,2051.8,1313.5,312.42,2773.3,1686.6,0.0000,6484.4,4449.7,4252.8,3658.0,0.0000,-362.55,-113.35,-77.419,-42.110,-96.171,-587.69,0.0000,-1076.3,-1599.9,-756.95,-1294.3
670.0000000000,91.676,1895.8,1960.6,1263.2,285.34,2591.0,972.43,1.7172,5386.5,2651.5,3352.4,1981.4,0.0000,-7347.4,-7185.9,-1597.9,-2583.3,-2859.9,-16879.,-155.89,-20315.,-6415.9,-4431.2,-2884.9,63.085,2247.4,2049.2,1309.5,311.99,2763.7,1686.6,0.0000,6478.6,4449.7,4252.8,3658.0,0.0000,-362.01,-113.16,-77.240,-42.057,-95.699,-587.69,0.0000,-1076.2,-1599.7,-756.94,-1294.1
671.0000000000,91.577,1893.4,1957.8,1259.1,284.88,2581.9,972.43,1.7177,5381.1,2651.6,3352.5,1981.6,0.0000,-7342.6,-7184.1,-1595.5,-2581.9,-2854.1,-16876.,-155.73,-20312.,-6415.5,-4430.5,-2883.9,63.006,2244.6,2046.7,1305.5,311.56,2754.2,1686.6,0.0000,6472.8,4449.7,4252.8,3658.0,0.0000,-361.48,-112.98,-77.063,-42.004,-95.229,-587.69,0.0000,-1076.1,-1599.5,-756.92,-1293.9
672.0000000000,91.482,1891.1,1955.3,1255.1,284.42,2572.7,972.43,1.7182,5375.4,2651.8,3352.5,1981.8,0.0000,-7337.9,-7182.3,-1593.1,-2580.6,-2848.3,-16873.,-155.56,-20309.,-6415.1,-4429.7,-2883.0,62.919,2241.5,2043.8,1301.3,311.09,2744.5,1686.6,0.0000,6466.9,4449.7,4252.8,3658.0,0.0000,-360.89,-112.78,-76.877,-41.946,-94.753,-587.69,0.0000,-1075.9,-1599.4,-756.90,-1293.7
673.0000000000,91.386,1888.7,1953.4,1251.2,284.01,2563.6,972.44,1.7188,5369.7,2651.9,3352.5,1982.0,0.0000,-7333.1,-7180.5,-1590.7,-2579.2,-2842.5,-16870.,-155.40,-20306.,-6414.6,-4429.0,-2882.0,62.821,2238.0,2040.7,1297.1,310.56,2734.4,1686.6,0.0000,6460.8,4449.7,4252.8,3658.0,0.0000,-360.24,-112.56,-76.679,-41.881,-94.266,-587.69,0.0000,-1075.8,-1599.2,-756.89,-1293.5
674.0000000000,91.317,1900.8,1964.7,1247.9,286.60,2556.3,972.44,1.7193,5364.2,2652.1,3352.5,1982.2,0.0000,-7329.6,-7179.3,-1588.6,-2577.9,-2836.8,-16867.,-155.24,-20303.,-6414.2,-4428.2,-2881.0,77.942,2367.6,2158.8,1338.0,328.46,2800.7,1686.6,81.162,6502.7,4455.1,4256.7,3663.3,0.0000,-378.12,-118.49,-79.589,-43.982,-96.417,-587.69,-3.7172,-1076.2,-1599.1,-756.89,-1293.6
675.0000000000,92.947,1948.2,2005.4,1250.8,294.22,2562.1,972.44,1.7198,5361.3,2652.2,3352.5,1982.3,0.0000,-7329.8,-7180.2,-1587.0,-2577.1,-2831.5,-16863.,-155.09,-20300.,-6413.8,-4427.4,-2880.1,719.34,3065.7,2874.0,1443.1,358.64,3017.0,1686.7,645.34,6642.0,4476.9,4274.9,3683.7,0.0000,-393.63,-136.54,-83.901,-45.773,-103.52,-587.69,-29.557,-1077.7,-1598.9,-756.97,-1294.2
676.0000000000,94.715,2002.4,2057.3,1269.4,301.62,2589.2,972.44,1.7204,5364.9,2652.4,3352.5,1982.5,0.0000,-7333.4,-7183.2,-1586.4,-2576.6,-2827.2,-16860.,-154.94,-20297.,-6413.4,-4426.7,-2879.1,69.959,2492.3,2272.5,1462.7,382.79,3033.2,1686.6,0.0000,6657.2,4474.3,4285.4,3697.8,0.0000,-401.10,-125.38,-85.000,-46.872,-103.76,-587.69,0.0000,-1077.8,-1598.7,-757.01,-1294.6
677.0000000000,96.322,2041.5,2096.7,1294.6,309.81,2619.9,972.44,1.7308,5371.5,2652.5,3352.5,1982.7,0.0000,-7338.9,-7186.9,-1585.9,-2576.3,-2823.9,-16857.,-154.78,-20294.,-6413.0,-4425.9,-2878.2,70.298,2504.3,2283.5,1445.0,358.18,3018.5,1686.6,0.0000,6636.5,4461.9,4264.1,3670.5,0.0000,-403.07,-126.03,-85.249,-46.934,-103.64,-587.69,0.0000,-1077.4,-1598.6,-756.88,-1293.3
678.0000000000,97.707,2061.6,2119.5,1313.3,313.88,2640.6,972.58,1.7322,5377.9,2652.7,3352.6,1982.9,0.0000,-7344.6,-7190.4,-1585.8,-2575.8,-2821.4,-16854.,-154.62,-20291.,-6412.5,-4425.1,-2877.2,70.398,2507.9,2286.8,1441.6,354.37,3014.9,1686.6,0.0000,6632.5,4457.2,4259.6,3665.4,0.0000,-403.69,-126.26,-85.316,-46.974,-103.54,-587.69,0.0000,-1077.3,-1598.4,-756.84,-1292.9
679.0000000000,98.462,2072.0,2132.0,1329.3,315.60,2653.4,972.59,1.7327,5381.3,2652.9,3352.5,1983.1,0.0000,-7349.7,-7193.5,-1585.6,-2575.3,-2818.4,-16851.,-154.46,-20289.,-6412.1,-4424.4,-2876.3,70.402,2508.0,2286.9,1438.1,350.87,3010.9,1686.6,0.0000,6628.6,4453.1,4255.9,3661.4,0.0000,-403.76,-126.32,-85.308,-46.954,-103.41,-587.69,0.0000,-1077.2,-1598.3,-756.80,-1292.5
680.0000000000,98.707,2077.9,2138.4,1338.0,315.90,2661.7,972.57,1.7332,5385.4,2653.0,3352.5,1983.3,0.0000,-7354.1,-7196.1,-1585.5,-2574.6,-2815.0,-16848.,-154.30,-20286.,-6411.7,-4423.6,-2875.3,70.349,2506.1,2285.2,1435.8,348.91,3007.8,1686.6,0.0000,6626.1,4451.2,4254.2,3659.5,0.0000,-403.50,-126.27,-85.251,-46.908,-103.27,-587.69,0.0000,-1077.1,-1598.1,-756.77,-1292.3
681.0000000000,98.727,2080.5,2143.9,1344.7,315.84,2665.3,972.55,2.2658,5392.9,2653.2,3352.6,1983.5,0.0000,-7357.9,-7198.3,-1585.6,-2573.9,-2811.4,-16845.,-154.14,-20283.,-6411.2,-4422.8,-2874.3,70.305,2504.6,2283.8,1434.5,347.86,3006.2,1686.6,0.0000,6624.8,4450.3,4253.4,3658.6,0.0000,-403.30,-126.24,-85.211,-46.874,-103.16,-587.69,0.0000,-1077.0,-1597.9,-756.75,-1292.0
682.0000000000,98.854,2083.7,2149.4,1346.9,315.64,2672.4,972.55,2.3143,5408.0,2653.2,3352.6,1983.7,0.0000,-7361.4,-7200.2,-1585.2,-2573.2,-2807.6,-16842.,-153.98,-20281.,-6410.8,-4422.1,-2873.4,70.255,2502.8,2282.1,1433.7,347.32,3005.1,1686.6,0.0000,6624.0,4450.0,4253.1,3658.3,0.0000,-403.05,-126.19,-85.167,-46.839,-103.05,-587.69,0.0000,-1076.9,-1597.8,-756.73,-1291.8
683.0000000000,98.837,2086.7,2152.3,1348.0,315.36,2691.1,972.53,2.3148,5429.3,2653.5,3352.6,1983.9,0.0000,-7364.6,-7201.8,-1584.6,-2572.3,-2803.6,-16839.,-153.82,-20278.,-6410.4,-4421.3,-2872.4,70.204,2501.0,2280.5,1433.0,346.93,3004.1,1686.6,0.0000,6623.3,4449.8,4252.9,3658.1,0.0000,-402.80,-126.13,-85.122,-46.804,-102.94,-587.69,0.0000,-1076.9,-1597.6,-756.71,-1291.6
684.0000000000,98.779,2087.3,2152.5,1349.5,315.09,2710.2,972.49,2.3153,5443.4,2653.6,3352.6,1984.1,0.0000,-7367.4,-7203.2,-1583.8,-2571.5,-2799.7,-16836.,-153.66,-20275.,-6410.0,-4420.5,-2871.5,70.132,2498.4,2278.1,1432.0,346.50,3002.3,1686.6,0.0000,6622.2,4449.7,4252.8,3658.0,0.0000,-402.41,-126.03,-85.051,-46.755,-102.81,-587.69,0.0000,-1076.8,-1597.5,-756.70,-1291.5
685.0000000000,98.709,2088.2,2151.3,1351.6,314.79,2721.2,972.49,2.3158,5450.6,2653.8,3352.7,1984.3,0.0000,-7369.5,-7204.3,-1582.9,-2570.7,-2795.7,-16832.,-153.51,-20273.,-6409.5,-4419.8,-2870.5,70.037,2495.0,2275.0,1430.5,346.00,2999.6,1686.6,0.0000,6620.6,4449.7,4252.8,3658.0,0.0000,-401.89,-125.89,-84.953,-46.691,-102.64,-587.69,0.0000,-1076.7,-1597.3,-756.68,-1291.3
686.0000000000,98.624,2089.4,2151.4,1353.1,314.44,2723.4,972.49,2.7592,5454.1,2654.0,3352.7,1984.5,0.0000,-7371.1,-7205.3,-1582.0,-2569.8,-2791.7,-16829.,-153.35,-20270.,-6409.1,-4419.0,-2869.5,69.955,2492.1,2272.4,1429.2,345.58,2997.2,1686.6,0.0000,6619.1,4449.7,4252.8,3658.0,0.0000,-401.45,-125.77,-84.868,-46.637,-102.47,-587.69,0.0000,-1076.6,-1597.2,-756.66,-1291.1
687.0000000000,98.538,2088.3,2151.4,1353.6,314.09,2722.4,972.49,3.6754,5455.3,2654.1,3352.7,1984.7,0.0000,-7372.3,-7206.2,-1581.0,-2568.9,-2787.7,-16826.,-153.19,-20268.,-6408.7,-4418.2,-2868.6,69.871,2489.1,2269.7,1427.7,345.16,2994.4,1686.6,0.0000,6617.5,4449.7,4252.8,3658.0,0.0000,-400.98,-125.64,-84.775,-46.581,-102.30,-587.69,0.0000,-1076.6,-1597.0,-756.64,-1290.9
688.0000000000,98.375,2087.4,2150.4,1352.8,313.72,2719.8,972.49,3.6758,5454.1,2654.2,3352.7,1984.9,0.0000,-7373.1,-7207.0,-1580.0,-2568.0,-2783.7,-16823.,-153.03,-20265.,-6408.2,-4417.5,-2867.6,69.776,2485.7,2266.6,1426.0,344.70,2991.0,1686.6,0.0000,6615.5,4449.7,4252.8,3658.0,0.0000,-400.45,-125.48,-84.668,-46.517,-102.11,-587.69,0.0000,-1076.5,-1596.9,-756.63,-1290.7
689.0000000000,98.256,2085.7,2151.0,1351.5,313.31,2718.4,972.49,4.1936,5452.7,2654.3,3352.7,1985.1,0.0000,-7373.8,-7207.6,-1578.9,-2567.1,-2779.7,-16820.,-152.88,-20263.,-6407.8,-4416.7,-2866.7,69.662,2481.7,2262.9,1423.9,344.14,2986.8,1686.6,0.0000,6612.9,4449.7,4252.8,3658.0,0.0000,-399.80,-125.29,-84.537,-46.441,-101.88,-587.69,0.0000,-1076.4,-1596.7,-756.61,-1290.5
690.0000000000,98.146,2083.5,2149.6,1350.0,312.85,2719.9,972.49,4.5946,5453.4,2654.5,3352.7,1985.3,0.0000,-7374.3,-7208.1,-1577.7,-2566.1,-2775.8,-16817.,-152.73,-20260.,-6407.4,-4415.9,-2865.7,69.533,2477.1,2258.7,1421.4,343.50,2981.9,1686.6,0.0000,6609.9,4449.7,4252.8,3658.0,0.0000,-399.06,-125.07,-84.386,-46.355,-101.63,-587.69,0.0000,-1076.3,-1596.5,-756.59,-1290.3
691.0000000000,98.023,2081.6,2146.4,1348.7,312.33,2719.4,972.49,5.6165,5454.3,2654.7,3352.7,1985.5,0.0000,-7374.4,-7208.4,-1576.6,-2565.1,-2771.9,-16814.,-152.57,-20258.,-6406.9,-4415.1,-2864.7,69.388,2471.9,2254.0,1418.6,342.79,2976.1,1686.6,0.0000,6606.4,4449.7,4252.8,3658.0,0.0000,-398.23,-124.82,-84.213,-46.258,-101.35,-587.69,0.0000,-1076.2,-1596.4,-756.57,-1290.1
692.0000000000,97.889,2079.4,2143.5,1348.3,311.94,2720.0,972.49,5.6167,5452.9,2654.8,3352.8,1985.7,0.0000,-7374.3,-7208.5,-1575.4,-2564.2,-2768.0,-16811.,-152.42,-20255.,-6406.5,-4414.4,-2863.8,69.460,2474.5,2312.1,1420.8,386.17,2981.1,1686.6,0.0000,6609.5,4449.7,4252.8,3658.0,0.0000,-398.64,-126.14,-84.328,-46.576,-101.45,-587.69,0.0000,-1076.2,-1596.2,-756.56,-1289.9
693.0000000000,97.860,2078.1,2141.9,1347.5,311.75,2718.8,972.50,5.6439,5451.1,2655.0,3352.8,1985.9,0.0000,-7374.1,-7208.6,-1574.2,-2563.2,-2764.1,-16808.,-152.28,-20253.,-6406.0,-4413.6,-2862.8,69.343,2470.3,2252.5,1418.2,342.57,2975.5,1686.6,0.0000,6606.1,4449.7,4252.8,3658.0,0.0000,-397.96,-124.75,-84.177,-46.228,-101.18,-587.69,0.0000,-1076.1,-1596.1,-756.54,-1289.8
694.0000000000,97.749,2075.8,2139.7,1346.7,311.38,2716.5,972.50,5.6999,5450.4,2655.2,3352.8,1986.1,0.0000,-7373.6,-7208.6,-1572.9,-2562.2,-2760.3,-16805.,-152.13,-20250.,-6405.6,-4412.8,-2861.9,69.246,2466.8,2249.4,1415.8,342.09,2970.5,1686.6,0.0000,6603.1,4449.7,4252.8,3658.0,0.0000,-397.39,-124.57,-84.046,-46.164,-100.93,-587.69,0.0000,-1076.0,-1595.9,-756.52,-1289.6
695.0000000000,97.645,2073.8,2136.9,1345.2,311.08,2713.2,972.54,5.7067,5450.6,2655.3,3352.9,1986.3,0.0000,-7372.9,-7208.4,-1571.7,-2561.2,-2756.4,-16802.,-151.98,-20248.,-6405.2,-4412.1,-2860.9,69.146,2463.3,2246.1,1413.4,341.59,2965.2,1686.6,0.0000,6599.9,4449.7,4252.8,3658.0,0.0000,-396.80,-124.39,-83.910,-46.097,-100.67,-587.69,0.0000,-1075.9,-1595.8,-756.51,-1289.4
696.0000000000,97.299,2071.7,2134.3,1344.4,310.62,2710.5,972.54,5.7069,5449.0,2655.5,3352.9,1986.4,0.0000,-7371.9,-7208.1,-1570.3,-2560.1,-2752.6,-16799.,-151.84,-20245.,-6404.7,-4411.3,-2859.9,69.032,2459.2,2242.4,1410.6,341.02,2959.3,1686.6,0.0000,6596.3,4449.7,4252.8,3658.0,0.0000,-396.13,-124.18,-83.757,-46.021,-100.39,-587.69,0.0000,-1075.8,-1595.6,-756.49,-1289.2
697.0000000000,97.183,2068.5,2131.9,1342.7,310.15,2708.0,972.54,5.7071,5448.3,2655.7,3352.9,1986.6,0.0000,-7370.8,-7207.6,-1569.0,-2559.1,-2748.7,-16796.,-151.70,-20243.,-6404.3,-4410.5,-2859.0,68.918,2455.2,2238.7,1407.8,340.45,2953.3,1686.6,0.0000,6592.7,4449.7,4252.8,3658.0,0.0000,-395.46,-123.97,-83.603,-45.946,-100.10,-587.69,0.0000,-1075.7,-1595.4,-756.47,-1289.0
698.0000000000,97.066,2065.5,2130.8,1340.8,309.66,2703.4,972.54,5.7074,5446.5,2655.8,3352.9,1986.8,0.0000,-7369.5,-7207.0,-1567.7,-2558.0,-2744.9,-16793.,-151.55,-20240.,-6403.9,-4409.8,-2858.0,68.799,2450.9,2234.8,1404.8,339.85,2946.9,1686.6,0.0000,6588.8,4449.7,4252.8,3658.0,0.0000,-394.75,-123.74,-83.439,-45.866,-99.805,-587.69,0.0000,-1075.6,-1595.3,-756.45,-1288.8
699.0000000000,96.943,2063.0,2129.9,1338.4,309.14,2701.0,972.54,7.3901,5444.4,2655.9,3352.9,1986.9,0.0000,-7368.1,-7206.3,-1566.3,-2557.0,-2741.0,-16790.,-151.41,-20238.,-6403.4,-4409.0,-2857.0,68.673,2446.4,2230.7,1401.6,339.22,2940.1,1686.6,0.0000,6584.7,4449.7,4252.8,3658.0,0.0000,-394.00,-123.50,-83.266,-45.782,-99.492,-587.69,0.0000,-1075.5,-1595.1,-756.44,-1288.6
700.0000000000,96.888,2059.9,2126.7,1335.8,308.61,2697.8,972.55,7.3158,5444.0,2656.0,3352.9,1987.1,0.0000,-7366.7,-7205.5,-1564.9,-2555.9,-2737.0,-16787.,-151.26,-20235.,-6403.0,-4408.2,-2856.1,68.548,2442.0,2226.7,1398.4,338.59,2933.2,1686.6,0.0000,6580.5,4449.7,4252.8,3658.0,0.0000,-393.25,-123.27,-83.093,-45.699,-99.177,-587.69,0.0000,-1075.4,-1595.0,-756.42,-1288.4
701.0000000000,96.859,2056.6,2123.5,1333.9,308.10,2693.1,972.55,5.6314,5445.7,2656.2,3353.0,1987.3,0.0000,-7365.0,-7204.6,-1563.4,-2554.8,-2733.0,-16785.,-151.12,-20233.,-6402.5,-4407.5,-2855.1,68.460,2438.8,2223.8,1395.8,338.14,2927.4,1686.6,0.0000,6577.0,4449.7,4252.8,3658.0,0.0000,-392.71,-123.09,-82.957,-45.640,-98.897,-587.69,0.0000,-1075.3,-1594.8,-756.40,-1288.3
702.0000000000,96.747,2053.7,2122.8,1331.7,307.64,2688.7,972.55,5.7039,5443.4,2656.4,3353.0,1987.5,0.0000,-7363.4,-7203.6,-1561.9,-2553.7,-2729.0,-16782.,-150.98,-20230.,-6402.1,-4406.7,-2854.1,68.360,2435.3,2220.6,1393.0,337.63,2921.1,1686.6,0.0000,6573.2,4449.7,4252.8,3658.0,0.0000,-392.10,-122.89,-82.808,-45.574,-98.600,-587.69,0.0000,-1075.2,-1594.7,-756.38,-1288.1
703.0000000000,96.603,2051.0,2120.8,1329.0,307.17,2685.4,972.55,7.5734,5441.1,2656.6,3353.0,1987.7,0.0000,-7361.6,-7202.6,-1560.4,-2552.6,-2724.9,-16779.,-150.84,-20228.,-6401.7,-4405.9,-2853.2,68.246,2431.2,2216.9,1389.8,337.05,2914.2,1686.6,0.0000,6569.0,4449.7,4252.8,3658.0,0.0000,-391.41,-122.67,-82.642,-45.497,-98.284,-587.69,0.0000,-1075.1,-1594.5,-756.37,-1287.9
704.0000000000,96.350,2047.4,2117.4,1326.3,306.71,2680.4,972.52,7.5735,5439.3,2656.7,3353.0,1987.9,0.0000,-7359.6,-7201.5,-1558.9,-2551.4,-2720.9,-16776.,-150.69,-20225.,-6401.2,-4405.2,-2852.2,68.124,2426.9,2212.9,1386.5,336.43,2906.9,1686.6,0.0000,6564.6,4449.7,4252.8,3658.0,0.0000,-390.67,-122.43,-82.464,-45.416,-97.953,-587.69,0.0000,-1074.9,-1594.4,-756.35,-1287.7
705.0000000000,96.358,2044.0,2113.9,1323.5,306.21,2676.1,972.51,7.5735,5436.1,2656.9,3353.0,1988.1,0.0000,-7357.5,-7200.3,-1557.3,-2550.3,-2716.9,-16773.,-150.55,-20222.,-6400.8,-4404.4,-2851.2,68.003,2422.6,2209.0,1383.1,335.82,2899.5,1686.6,0.0000,6560.1,4449.7,4252.8,3658.0,0.0000,-389.93,-122.19,-82.287,-45.335,-97.619,-587.69,0.0000,-1074.8,-1594.2,-756.33,-1287.5
706.0000000000,96.271,2040.6,2110.5,1320.5,305.69,2671.0,972.51,6.3692,5432.7,2657.0,3353.0,1988.2,0.0000,-7355.3,-7199.1,-1555.7,-2549.1,-2712.9,-16770.,-150.41,-20220.,-6400.3,-4403.6,-2850.3,67.889,2418.5,2205.3,1379.8,335.24,2892.1,1686.6,0.0000,6555.7,4449.7,4252.8,3658.0,0.0000,-389.23,-121.96,-82.114,-45.259,-97.287,-587.69,0.0000,-1074.7,-1594.1,-756.31,-1287.3
707.0000000000,96.096,2037.3,2107.1,1317.5,305.18,2666.1,972.51,5.5541,5429.3,2657.2,3353.1,1988.4,0.0000,-7352.8,-7197.8,-1554.1,-2548.0,-2708.8,-16767.,-150.27,-20217.,-6399.9,-4402.9,-2849.3,67.781,2414.7,2201.8,1376.5,334.69,2884.9,1686.6,0.0000,6551.3,4449.7,4252.8,3658.0,0.0000,-388.56,-121.74,-81.948,-45.187,-96.959,-587.69,0.0000,-1074.6,-1593.9,-756.30,-1287.1
708.0000000000,95.868,2034.1,2103.7,1314.4,304.71,2660.0,972.51,5.5542,5425.8,2657.3,3353.1,1988.6,0.0000,-7350.2,-7196.5,-1552.5,-2546.8,-2704.7,-16764.,-150.13,-20215.,-6399.5,-4402.1,-2848.3,67.671,2410.8,2198.2,1373.2,334.13,2877.6,1686.6,0.0000,6546.9,4449.7,4252.8,3658.0,0.0000,-387.89,-121.52,-81.779,-45.114,-96.627,-587.69,0.0000,-1074.5,-1593.8,-756.28,-1287.0
709.0000000000,95.749,2030.9,2100.5,1311.3,304.22,2655.5,972.50,5.5544,5422.2,2657.5,3353.1,1988.8,0.0000,-7347.5,-7195.1,-1550.8,-2545.7,-2700.6,-16761.,-149.98,-20212.,-6399.0,-4401.3,-2847.4,67.560,2406.8,2194.6,1369.8,333.56,2870.0,1686.6,0.0000,6542.3,4449.7,4252.8,3658.0,0.0000,-387.20,-121.29,-81.605,-45.040,-96.288,-587.69,0.0000,-1074.4,-1593.6,-756.26,-1286.8
710.0000000000,95.632,2027.7,2097.5,1308.2,303.74,2649.7,972.45,5.5545,5418.5,2657.6,3353.1,1989.0,0.0000,-7344.7,-7193.7,-1549.2,-2544.5,-2696.4,-16758.,-149.84,-20210.,-6398.6,-4400.6,-2846.4,67.467,2403.5,2191.6,1366.6,333.08,2862.7,1686.6,0.0000,6537.8,4449.7,4252.8,3658.0,0.0000,-386.61,-121.09,-81.447,-44.978,-95.955,-587.69,0.0000,-1074.3,-1593.4,-756.24,-1286.6
711.0000000000,95.524,2024.8,2094.4,1305.1,303.29,2643.7,972.43,5.5547,5414.8,2657.8,3353.1,1989.2,0.0000,-7341.8,-7192.3,-1547.5,-2543.3,-2692.1,-16755.,-149.70,-20207.,-6398.1,-4399.8,-2845.4,67.354,2399.4,2187.9,1363.1,332.50,2855.0,1686.6,0.0000,6533.2,4449.7,4252.8,3658.0,0.0000,-385.91,-120.86,-81.270,-44.902,-95.610,-587.69,0.0000,-1074.2,-1593.3,-756.23,-1286.4
712.0000000000,95.423,2021.5,2091.3,1302.0,302.79,2638.8,972.43,6.0552,5411.7,2658.0,3353.1,1989.4,0.0000,-7338.8,-7190.9,-1545.8,-2542.1,-2687.9,-16752.,-149.56,-20205.,-6397.7,-4399.0,-2844.5,67.237,2395.3,2184.1,1359.6,331.90,2847.1,1686.6,0.0000,6528.4,4449.7,4252.8,3658.0,0.0000,-385.18,-120.62,-81.089,-44.825,-95.259,-587.69,0.0000,-1074.1,-1593.1,-756.21,-1286.2
713.0000000000,95.481,2018.2,2087.9,1298.8,302.30,2632.3,972.39,7.5015,5409.0,2658.2,3353.2,1989.6,0.0000,-7335.7,-7189.4,-1544.1,-2540.9,-2683.6,-16750.,-149.42,-20202.,-6397.2,-4398.3,-2843.5,67.121,2391.1,2180.3,1356.0,331.31,2839.2,1686.6,0.0000,6523.6,4449.7,4252.8,3658.0,0.0000,-384.46,-120.38,-80.908,-44.747,-94.907,-587.69,0.0000,-1074.0,-1593.0,-756.19,-1286.0
714.0000000000,95.361,2014.9,2084.2,1295.6,301.79,2626.0,972.39,7.5015,5405.1,2658.4,3353.2,1989.8,0.0000,-7332.4,-7187.8,-1542.3,-2539.7,-2679.2,-16747.,-149.28,-20200.,-6396.8,-4397.5,-2842.6,67.012,2387.3,2176.8,1352.6,330.75,2831.4,1686.6,0.0000,6518.9,4449.7,4252.8,3658.0,0.0000,-383.77,-120.15,-80.733,-44.675,-94.561,-587.69,0.0000,-1073.8,-1592.8,-756.17,-1285.8
715.0000000000,95.242,2011.6,2080.8,1292.3,301.30,2620.7,972.39,7.0785,5402.0,2658.5,3353.2,1990.0,0.0000,-7329.1,-7186.3,-1540.6,-2538.5,-2674.9,-16744.,-149.14,-20197.,-6396.4,-4396.8,-2841.6,66.907,2383.5,2173.4,1349.2,330.21,2823.7,1686.6,0.0000,6514.3,4449.7,4252.8,3658.0,0.0000,-383.11,-119.93,-80.562,-44.605,-94.216,-587.69,0.0000,-1073.7,-1592.7,-756.16,-1285.7
716.0000000000,95.126,2008.6,2077.6,1289.1,300.82,2614.1,972.39,5.4794,5398.1,2658.7,3353.3,1990.2,0.0000,-7325.7,-7184.7,-1538.8,-2537.3,-2670.5,-16741.,-149.00,-20195.,-6395.9,-4396.0,-2840.6,66.815,2380.2,2170.4,1345.9,329.73,2816.4,1686.6,0.0000,6509.8,4449.7,4252.8,3658.0,0.0000,-382.52,-119.73,-80.405,-44.543,-93.884,-587.69,0.0000,-1073.6,-1592.5,-756.14,-1285.5
717.0000000000,95.019,2005.6,2074.6,1285.8,300.38,2607.4,972.40,5.4795,5394.2,2658.9,3353.3,1990.3,0.0000,-7322.3,-7183.1,-1537.0,-2536.1,-2666.1,-16738.,-148.86,-20192.,-6395.5,-4395.2,-2839.7,66.722,2376.9,2167.4,1342.7,329.25,2809.0,1686.6,0.0000,6505.4,4449.7,4252.8,3658.0,0.0000,-381.93,-119.53,-80.246,-44.481,-93.550,-587.69,0.0000,-1073.5,-1592.4,-756.12,-1285.3
718.0000000000,94.914,2002.9,2071.8,1282.6,299.98,2600.7,972.40,5.4796,5390.3,2659.1,3353.3,1990.5,0.0000,-7318.8,-7181.5,-1535.3,-2534.9,-2661.7,-16735.,-148.72,-20190.,-6395.0,-4394.5,-2838.7,66.654,2374.5,2165.2,1339.6,328.89,2801.8,1686.6,0.0000,6501.0,4449.7,4252.8,3658.0,0.0000,-381.47,-119.38,-80.106,-44.436,-93.222,-587.69,0.0000,-1073.4,-1592.2,-756.10,-1285.1
719.0000000000,94.826,2000.4,2069.1,1279.5,299.61,2594.2,972.40,5.1885,5388.0,2659.3,3353.3,1990.7,0.0000,-7315.3,-7179.9,-1533.5,-2533.7,-2657.3,-16732.,-148.58,-20187.,-6394.6,-4393.7,-2837.7,66.565,2371.4,2162.3,1336.4,328.42,2794.5,1686.6,0.0000,6496.6,4449.7,4252.8,3658.0,0.0000,-380.90,-119.18,-79.951,-44.377,-92.891,-587.69,0.0000,-1073.3,-1592.1,-756.09,-1284.9
720.0000000000,94.732,1998.1,2066.4,1276.4,299.20,2587.5,972.40,3.4684,5384.4,2659.7,3353.3,1990.9,0.0000,-7311.7,-7178.2,-1531.7,-2532.4,-2652.9,-16729.,-148.44,-20184.,-6394.1,-4392.9,-2836.8,66.476,2368.2,2159.4,1333.2,327.96,2787.1,1686.6,0.0000,6492.1,4449.7,4252.8,3658.0,0.0000,-380.33,-118.99,-79.795,-44.317,-92.559,-587.69,0.0000,-1073.2,-1591.9,-756.07,-1284.7
721.0000000000,94.639,1996.4,2063.6,1273.3,298.82,2580.9,972.40,3.4739,5380.9,2659.9,3353.4,1991.1,0.0000,-7308.1,-7176.6,-1529.9,-2531.2,-2648.4,-16726.,-148.30,-20182.,-6393.7,-4392.2,-2835.8,66.388,2365.0,2156.5,1330.0,327.50,2779.8,1686.6,0.0000,6487.7,4449.7,4252.8,3658.0,0.0000,-379.76,-118.79,-79.640,-44.259,-92.227,-587.69,0.0000,-1073.1,-1591.8,-756.05,-1284.6
722.0000000000,94.546,1993.8,2061.0,1270.2,298.43,2574.1,972.40,3.4741,5376.9,2660.1,3353.4,1991.3,0.0000,-7304.5,-7175.0,-1528.0,-2530.0,-2644.0,-16723.,-148.17,-20179.,-6393.3,-4391.4,-2834.9,66.310,2362.3,2154.0,1326.9,327.09,2772.5,1686.6,0.0000,6483.2,4449.7,4252.8,3658.0,0.0000,-379.25,-118.62,-79.492,-44.207,-91.895,-587.69,0.0000,-1073.0,-1591.6,-756.03,-1284.4
723.0000000000,94.457,1991.6,2058.6,1267.1,298.09,2567.5,972.35,3.4744,5372.9,2660.2,3353.4,1991.5,0.0000,-7300.8,-7173.4,-1526.2,-2528.8,-2639.5,-16721.,-148.03,-20177.,-6392.8,-4390.7,-2833.9,66.270,2360.8,2152.7,1324.4,326.86,2766.5,1686.6,0.0000,6479.6,4449.7,4252.8,3658.0,0.0000,-378.95,-118.51,-79.386,-44.180,-91.610,-587.69,0.0000,-1072.9,-1591.5,-756.02,-1284.2
724.0000000000,94.388,1989.8,2056.5,1264.9,297.79,2561.0,972.26,3.4746,5369.0,2660.4,3353.4,1991.6,0.0000,-7297.2,-7171.8,-1524.4,-2527.6,-2635.0,-16718.,-147.89,-20174.,-6392.4,-4389.9,-2833.0,66.197,2358.2,2150.3,1321.4,326.48,2759.6,1686.6,0.0000,6475.4,4449.7,4252.8,3658.0,0.0000,-378.46,-118.34,-79.247,-44.131,-91.292,-587.69,0.0000,-1072.8,-1591.3,-756.00,-1284.0
725.0000000000,94.383,1987.7,2054.0,1262.2,297.46,2554.6,972.18,3.4749,5365.1,2660.5,3353.4,1991.8,0.0000,-7293.6,-7170.1,-1522.6,-2526.3,-2630.5,-16715.,-147.75,-20171.,-6391.9,-4389.1,-2832.0,66.110,2355.1,2147.5,1318.2,326.02,2752.2,1686.6,0.0000,6471.0,4449.7,4252.8,3658.0,0.0000,-377.90,-118.15,-79.092,-44.074,-90.959,-587.69,0.0000,-1072.7,-1591.2,-755.98,-1283.8
726.0000000000,94.419,1985.4,2051.4,1259.3,297.12,2548.2,972.17,3.4752,5361.2,2660.7,3353.4,1992.0,0.0000,-7289.9,-7168.5,-1520.7,-2525.1,-2626.0,-16712.,-147.61,-20169.,-6391.5,-4388.4,-2831.0,66.012,2351.7,2144.3,1314.8,325.52,2744.4,1686.6,0.0000,6466.3,4449.7,4252.8,3658.0,0.0000,-377.27,-117.94,-78.925,-44.008,-90.614,-587.69,0.0000,-1072.6,-1591.0,-755.96,-1283.6
727.0000000000,94.340,1986.3,2052.2,1256.7,297.36,2542.6,972.17,3.4786,5357.4,2660.8,3353.5,1992.2,0.0000,-7286.5,-7167.0,-1519.0,-2523.9,-2621.5,-16709.,-147.48,-20166.,-6391.1,-4387.6,-2830.1,70.356,2386.1,2181.2,1330.2,332.61,2774.1,1686.6,3.6684,6484.8,4451.3,4254.6,3660.0,0.0000,-381.12,-119.44,-79.744,-44.486,-91.487,-587.69,-0.16798,-1072.7,-1590.9,-755.96,-1283.5
728.0000000000,94.655,1994.3,2058.7,1255.9,298.59,2540.2,972.15,3.4768,5354.5,2661.0,3353.5,1992.4,0.0000,-7283.8,-7165.9,-1517.3,-2522.8,-2617.1,-16706.,-147.34,-20164.,-6390.6,-4386.9,-2829.1,66.912,2383.7,2173.6,1328.3,329.95,2769.5,1686.6,0.0000,6481.3,4449.7,4252.8,3658.0,0.0000,-382.30,-119.49,-79.851,-44.609,-91.300,-587.69,0.0000,-1072.6,-1590.7,-755.93,-1283.3
729.0000000000,94.822,2000.0,2064.5,1257.6,299.27,2538.8,972.13,3.4771,5352.0,2661.2,3353.5,1992.6,0.0000,-7281.5,-7165.1,-1515.7,-2521.7,-2612.8,-16703.,-147.21,-20161.,-6390.2,-4386.1,-2828.2,66.921,2384.0,2173.8,1325.9,329.94,2763.2,1686.6,0.0000,6477.5,4449.7,4252.8,3658.0,0.0000,-382.30,-119.48,-79.774,-44.614,-91.006,-587.69,0.0000,-1072.5,-1590.6,-755.91,-1283.1
730.0000000000,94.963,2002.4,2067.0,1258.2,300.02,2536.7,972.13,1.8200,5349.6,2661.3,3353.5,1992.7,0.0000,-7279.3,-7164.3,-1514.2,-2520.6,-2608.7,-16700.,-147.07,-20158.,-6389.7,-4385.3,-2827.2,66.944,2384.9,2174.6,1324.2,330.02,2758.4,1686.6,0.0000,6474.5,4449.7,4252.8,3658.0,0.0000,-382.38,-119.50,-79.726,-44.630,-90.762,-587.69,0.0000,-1072.4,-1590.4,-755.89,-1282.9
731.0000000000,95.113,2004.1,2068.8,1258.2,300.37,2533.6,972.13,1.4516,5347.1,2661.5,3353.5,1992.9,0.0000,-7277.2,-7163.5,-1512.6,-2519.6,-2604.5,-16698.,-146.94,-20156.,-6389.3,-4384.6,-2826.3,67.067,2389.2,2178.6,1324.3,330.57,2757.2,1686.6,0.0000,6473.8,4449.7,4252.8,3658.0,0.0000,-383.03,-119.70,-79.792,-44.712,-90.642,-587.69,0.0000,-1072.3,-1590.3,-755.88,-1282.7
732.0000000000,95.205,2007.1,2071.4,1257.7,300.75,2530.3,972.11,1.4522,5344.3,2661.6,3353.5,1993.1,0.0000,-7275.2,-7162.8,-1511.1,-2518.5,-2600.2,-16695.,-146.80,-20153.,-6388.9,-4383.8,-2825.3,69.695,2415.2,2195.8,1331.4,332.56,2761.2,1686.6,2.8902,6479.0,4451.1,4253.1,3658.0,0.0000,-384.14,-120.26,-79.938,-44.849,-90.618,-587.69,-0.13234,-1072.3,-1590.1,-755.86,-1282.6
733.0000000000,95.222,2011.7,2075.5,1257.5,301.39,2528.3,972.11,1.4527,5342.5,2661.5,3353.5,1993.3,0.0000,-7273.5,-7162.2,-1509.6,-2517.4,-2596.0,-16692.,-146.67,-20150.,-6388.4,-4383.1,-2824.4,77.844,2440.3,2234.4,1339.5,343.08,2771.7,1686.6,7.9873,6486.8,4456.6,4261.7,3665.8,0.0000,-385.62,-121.35,-80.143,-45.082,-90.660,-587.69,-0.36573,-1072.4,-1590.0,-755.89,-1282.7
734.0000000000,95.576,2016.5,2080.5,1257.7,302.12,2525.9,972.11,1.4532,5340.9,2661.6,3353.5,1993.4,0.0000,-7272.1,-7161.8,-1508.2,-2516.4,-2591.8,-16689.,-146.53,-20148.,-6388.0,-4382.3,-2823.4,67.597,2408.1,2195.8,1325.8,333.00,2755.2,1686.6,0.0000,6472.5,4449.7,4252.8,3658.0,0.0000,-385.94,-120.60,-80.116,-45.065,-90.335,-587.69,0.0000,-1072.1,-1589.8,-755.82,-1282.2
735.0000000000,95.720,2020.0,2084.3,1257.5,302.58,2524.3,972.11,1.4537,5341.2,2661.7,3353.5,1993.6,0.0000,-7270.8,-7161.4,-1506.7,-2515.4,-2587.6,-16686.,-146.40,-20145.,-6387.5,-4381.5,-2822.5,67.616,2408.8,2196.4,1323.6,333.05,2749.2,1686.6,0.0000,6468.8,4449.7,4252.8,3658.0,0.0000,-386.01,-120.61,-80.049,-45.077,-90.053,-587.69,0.0000,-1072.0,-1589.7,-755.81,-1282.0
736.0000000000,95.811,2021.6,2085.9,1256.9,302.85,2523.2,972.11,1.4543,5340.7,2661.9,3353.5,1993.8,0.0000,-7269.4,-7161.0,-1505.2,-2514.4,-2583.5,-16683.,-146.26,-20142.,-6387.1,-4380.8,-2821.5,67.600,2408.2,2195.9,1321.0,332.93,2742.8,1686.6,0.0000,6464.9,4449.7,4252.8,3658.0,0.0000,-385.88,-120.57,-79.954,-45.067,-89.759,-587.69,0.0000,-1071.9,-1589.5,-755.79,-1281.8
737.0000000000,95.939,2021.8,2086.2,1255.9,302.82,2521.1,972.08,1.4598,5339.5,2662.1,3353.5,1994.0,0.0000,-7268.0,-7160.5,-1503.7,-2513.3,-2579.2,-16680.,-146.13,-20140.,-6386.7,-4380.0,-2820.6,67.547,2406.3,2194.2,1318.0,332.63,2735.6,1686.6,0.0000,6460.6,4449.7,4252.8,3658.0,0.0000,-385.54,-120.46,-79.825,-45.031,-89.440,-587.69,0.0000,-1071.8,-1589.4,-755.77,-1281.7
738.0000000000,96.011,2021.8,2085.9,1254.5,302.67,2517.1,972.08,1.4687,5337.7,2662.2,3353.5,1994.2,0.0000,-7266.4,-7159.9,-1502.2,-2512.3,-2574.9,-16678.,-145.99,-20137.,-6386.2,-4379.3,-2819.6,67.509,2405.0,2192.9,1315.4,332.40,2729.2,1686.6,0.0000,6456.7,4449.7,4252.8,3658.0,0.0000,-385.29,-120.38,-79.715,-45.006,-89.146,-587.69,0.0000,-1071.7,-1589.2,-755.75,-1281.5
739.0000000000,95.976,2021.5,2085.8,1252.6,302.49,2512.5,972.08,1.4693,5335.8,2662.3,3353.6,1994.4,0.0000,-7264.6,-7159.3,-1500.6,-2511.2,-2570.6,-16675.,-145.86,-20135.,-6385.8,-4378.5,-2818.7,67.478,2403.9,2191.9,1313.1,332.22,2723.5,1686.6,0.0000,6453.2,4449.7,4252.8,3658.0,0.0000,-385.08,-120.31,-79.620,-44.985,-88.876,-587.69,0.0000,-1071.6,-1589.1,-755.74,-1281.3
740.0000000000,95.779,2022.8,2087.3,1250.7,302.64,2508.2,972.08,1.4698,5334.6,2662.4,3353.6,1994.5,0.0000,-7263.0,-7158.7,-1499.1,-2510.1,-2566.3,-16672.,-145.72,-20132.,-6385.3,-4377.7,-2817.7,76.630,2461.7,2242.8,1333.4,343.33,2744.9,1686.6,0.24049,6467.5,4451.6,4263.1,3665.2,0.0000,-387.25,-121.79,-79.955,-45.292,-89.098,-587.69,-0.11011E-01,-1071.7,-1588.9,-755.77,-1281.4
741.0000000000,95.948,2027.8,2091.3,1249.2,303.28,2505.4,972.08,1.4703,5333.1,2662.5,3353.6,1994.7,0.0000,-7261.7,-7158.3,-1497.5,-2509.1,-2562.0,-16669.,-145.59,-20129.,-6384.9,-4377.0,-2816.8,67.921,2419.6,2206.3,1315.9,334.29,2725.7,1686.6,0.0000,6454.5,4449.7,4252.8,3658.0,0.0000,-387.54,-121.07,-79.942,-45.281,-88.793,-587.69,0.0000,-1071.5,-1588.8,-755.70,-1281.0
742.0000000000,96.013,2030.6,2094.3,1249.3,303.55,2503.2,972.08,1.4708,5331.2,2662.6,3353.7,1994.9,0.0000,-7260.6,-7158.0,-1496.0,-2508.1,-2557.8,-16666.,-145.45,-20127.,-6384.4,-4376.2,-2815.8,67.894,2418.7,2205.4,1313.2,334.13,2719.2,1686.6,0.0000,6450.5,4449.7,4252.8,3658.0,0.0000,-387.35,-121.02,-79.838,-45.263,-88.496,-587.69,0.0000,-1071.4,-1588.6,-755.68,-1280.8
743.0000000000,96.072,2031.6,2095.0,1248.5,303.83,2500.4,972.08,1.4713,5329.1,2662.8,3353.6,1995.0,0.0000,-7259.3,-7157.7,-1494.4,-2507.1,-2553.6,-16663.,-145.32,-20124.,-6384.0,-4375.5,-2814.9,67.850,2417.1,2204.0,1310.5,333.88,2712.5,1686.6,0.0000,6446.5,4449.7,4252.8,3658.0,0.0000,-387.07,-120.92,-79.721,-45.233,-88.194,-587.69,0.0000,-1071.3,-1588.5,-755.67,-1280.6
744.0000000000,96.101,2031.4,2094.9,1247.3,303.74,2496.3,972.08,1.4770,5326.5,2663.0,3353.7,1995.2,0.0000,-7257.9,-7157.2,-1492.9,-2506.1,-2549.4,-16660.,-145.19,-20122.,-6383.5,-4374.7,-2813.9,67.808,2415.6,2202.7,1307.9,333.64,2706.2,1686.6,0.0000,6442.7,4449.7,4252.8,3658.0,0.0000,-386.80,-120.84,-79.611,-45.206,-87.908,-587.69,0.0000,-1071.2,-1588.4,-755.65,-1280.4
745.0000000000,96.069,2030.7,2094.3,1245.7,303.53,2491.5,972.08,1.4904,5323.4,2663.1,3353.7,1995.4,0.0000,-7256.4,-7156.7,-1491.3,-2505.1,-2545.1,-16658.,-145.05,-20119.,-6383.1,-4373.9,-2813.0,67.754,2413.7,2200.9,1305.1,333.34,2699.7,1686.6,0.0000,6438.7,4449.7,4252.8,3658.0,0.0000,-386.46,-120.73,-79.489,-45.169,-87.614,-587.69,0.0000,-1071.1,-1588.2,-755.63,-1280.2
746.0000000000,96.014,2029.6,2093.4,1243.8,303.27,2486.5,972.08,1.5020,5320.4,2663.2,3353.7,1995.6,0.0000,-7254.7,-7156.1,-1489.7,-2504.0,-2540.9,-16655.,-144.92,-20116.,-6382.6,-4373.2,-2812.0,67.681,2411.1,2198.5,1302.2,332.96,2692.9,1686.6,0.0000,6434.6,4449.7,4252.8,3658.0,0.0000,-386.01,-120.58,-79.351,-45.121,-87.307,-587.69,0.0000,-1071.0,-1588.1,-755.61,-1280.1
747.0000000000,95.946,2028.1,2092.3,1241.5,302.95,2481.0,972.08,1.5025,5317.6,2663.4,3353.7,1995.7,0.0000,-7252.9,-7155.5,-1488.1,-2503.0,-2536.6,-16652.,-144.79,-20114.,-6382.2,-4372.4,-2811.1,67.596,2408.1,2195.8,1299.0,332.52,2685.7,1686.6,0.0000,6430.2,4449.7,4252.8,3658.0,0.0000,-385.49,-120.42,-79.200,-45.064,-86.992,-587.69,0.0000,-1070.9,-1587.9,-755.59,-1279.9
748.0000000000,95.867,2026.6,2090.7,1239.0,302.53,2476.0,972.09,1.5030,5315.6,2663.5,3353.7,1995.9,0.0000,-7251.0,-7154.7,-1486.5,-2501.9,-2532.3,-16649.,-144.65,-20111.,-6381.7,-4371.7,-2810.1,67.499,2404.6,2192.6,1295.7,332.01,2678.2,1686.6,0.0000,6425.7,4449.7,4252.8,3658.0,0.0000,-384.90,-120.23,-79.037,-44.999,-86.666,-587.69,0.0000,-1070.8,-1587.8,-755.58,-1279.7
749.0000000000,95.775,2024.4,2088.4,1236.6,302.12,2472.2,972.09,1.5035,5313.2,2663.7,3353.7,1996.0,0.0000,-7249.0,-7153.9,-1484.8,-2500.8,-2527.9,-16646.,-144.52,-20109.,-6381.3,-4370.9,-2809.2,67.400,2401.1,2189.4,1292.5,331.50,2670.8,1686.6,0.0000,6421.2,4449.7,4252.8,3658.0,0.0000,-384.29,-120.03,-78.873,-44.934,-86.341,-587.69,0.0000,-1070.7,-1587.6,-755.56,-1279.5
750.0000000000,95.675,2021.9,2086.0,1234.0,301.65,2467.5,972.09,1.5040,5310.5,2663.8,3353.7,1996.2,0.0000,-7246.8,-7153.0,-1483.1,-2499.7,-2523.6,-16643.,-144.39,-20106.,-6380.8,-4370.2,-2808.3,67.287,2397.1,2185.7,1288.9,330.92,2662.9,1686.6,0.0000,6416.4,4449.7,4252.8,3658.0,0.0000,-383.60,-119.81,-78.695,-44.858,-86.002,-587.69,0.0000,-1070.5,-1587.5,-755.54,-1279.4
751.0000000000,95.564,2019.3,2083.6,1231.3,301.18,2461.7,972.09,1.5045,5307.3,2664.0,3353.8,1996.4,0.0000,-7244.4,-7152.0,-1481.4,-2498.6,-2519.3,-16641.,-144.25,-20103.,-6380.4,-4369.4,-2807.3,67.169,2392.9,2181.9,1285.4,330.32,2655.0,1686.6,0.0000,6411.6,4449.7,4252.8,3658.0,0.0000,-382.89,-119.58,-78.512,-44.779,-85.661,-587.69,0.0000,-1070.4,-1587.3,-755.52,-1279.2
752.0000000000,95.449,2017.2,2081.7,1228.5,300.83,2455.8,972.09,1.5050,5303.8,2664.1,3353.8,1996.6,0.0000,-7242.0,-7151.0,-1479.7,-2497.5,-2514.9,-16638.,-144.12,-20101.,-6379.9,-4368.6,-2806.4,67.252,2395.8,2184.6,1285.2,330.70,2653.6,1686.6,1.8315,6413.1,4451.4,4252.8,3658.0,0.0000,-383.32,-119.70,-78.548,-44.835,-85.536,-587.69,-0.83854E-01,-1070.4,-1587.2,-755.51,-1279.0
753.0000000000,95.438,2017.9,2082.0,1226.0,300.91,2450.6,972.09,1.5055,5300.5,2664.2,3353.8,1996.8,0.0000,-7239.7,-7150.1,-1477.9,-2496.4,-2510.5,-16635.,-143.99,-20098.,-6379.5,-4367.9,-2805.4,70.681,2416.4,2199.2,1294.4,334.95,2660.7,1686.6,5.0594,6419.8,4455.0,4259.0,3663.4,0.0000,-384.25,-120.18,-78.678,-44.968,-85.536,-587.69,-0.23164,-1070.4,-1587.0,-755.52,-1279.0
754.0000000000,95.492,2019.7,2083.7,1224.3,301.09,2446.7,972.09,1.5060,5297.7,2664.3,3353.8,1996.9,0.0000,-7237.6,-7149.3,-1476.3,-2495.4,-2506.2,-16632.,-143.86,-20095.,-6379.0,-4367.1,-2804.5,67.392,2400.8,2189.1,1284.2,331.32,2649.3,1686.6,0.0000,6408.1,4449.7,4252.8,3658.0,0.0000,-384.03,-119.91,-78.585,-44.928,-85.241,-587.69,0.0000,-1070.2,-1586.9,-755.47,-1278.7
755.0000000000,95.491,2019.7,2084.1,1222.8,301.13,2442.4,972.09,1.5065,5294.6,2664.4,3353.9,1997.1,0.0000,-7235.6,-7148.5,-1474.6,-2494.3,-2501.9,-16629.,-143.73,-20093.,-6378.6,-4366.4,-2803.5,67.315,2398.1,2186.6,1281.2,330.92,2642.5,1686.6,0.0000,6404.0,4449.7,4252.8,3658.0,0.0000,-383.55,-119.75,-78.444,-44.877,-84.939,-587.69,0.0000,-1070.1,-1586.8,-755.45,-1278.5
756.0000000000,95.484,2018.5,2082.8,1221.0,301.06,2438.0,972.09,1.5070,5291.5,2664.5,3353.9,1973.9,0.0000,-7233.4,-7147.6,-1472.9,-2493.2,-2497.6,-16627.,-143.60,-20090.,-6378.1,-4365.6,-2802.6,67.222,2394.7,2183.6,1278.0,330.44,2635.3,1686.6,0.0000,6399.6,4449.7,4252.8,3658.0,0.0000,-382.97,-119.57,-78.287,-44.814,-84.623,-587.69,0.0000,-1070.0,-1586.6,-755.43,-1278.3
757.0000000000,95.433,2016.4,2081.0,1219.0,300.71,2432.8,972.09,1.5075,5288.4,2664.7,3353.9,1974.1,0.0000,-7231.2,-7146.7,-1471.2,-2492.2,-2493.4,-16624.,-143.47,-20088.,-6377.7,-4364.8,-2801.6,67.121,2391.2,2180.3,1274.7,329.92,2627.9,1686.6,0.0000,6395.2,4449.7,4252.8,3658.0,0.0000,-382.36,-119.37,-78.124,-44.748,-84.302,-587.69,0.0000,-1069.9,-1586.5,-755.42,-1278.1
758.0000000000,95.341,2013.8,2078.6,1216.8,300.28,2427.4,972.10,1.5080,5285.0,2664.8,3353.9,1974.3,0.0000,-7228.7,-7145.6,-1469.5,-2491.1,-2489.1,-16621.,-143.33,-20085.,-6377.2,-4364.1,-2800.7,67.003,2387.0,2176.5,1271.2,329.32,2620.0,1686.6,0.0000,6390.4,4449.7,4252.8,3658.0,0.0000,-381.64,-119.13,-77.942,-44.669,-83.966,-587.69,0.0000,-1069.8,-1586.3,-755.40,-1277.9
759.0000000000,95.229,2010.9,2075.7,1214.3,299.78,2421.4,972.10,1.5085,5281.6,2665.0,3353.9,1974.5,0.0000,-7226.2,-7144.5,-1467.8,-2489.9,-2484.7,-16618.,-143.20,-20082.,-6376.7,-4363.3,-2799.7,66.877,2382.4,2172.4,1267.5,328.67,2612.0,1686.6,0.0000,6385.5,4449.7,4252.8,3658.0,0.0000,-380.87,-118.88,-77.751,-44.584,-83.623,-587.69,0.0000,-1069.7,-1586.2,-755.38,-1277.8
760.0000000000,95.106,2007.9,2072.7,1211.5,299.26,2415.5,972.09,1.5090,5278.5,2665.1,3354.0,1974.7,0.0000,-7223.4,-7143.3,-1466.1,-2488.8,-2480.4,-16615.,-143.07,-20080.,-6376.3,-4362.6,-2798.8,66.751,2378.0,2168.3,1263.9,328.04,2604.0,1686.6,0.0000,6380.7,4449.7,4252.8,3658.0,0.0000,-380.12,-118.63,-77.563,-44.501,-83.283,-587.69,0.0000,-1069.6,-1586.0,-755.36,-1277.6
761.0000000000,94.981,2005.5,2070.3,1208.5,298.84,2409.8,972.09,1.5094,5275.8,2665.3,3354.0,1974.9,0.0000,-7220.7,-7142.1,-1464.3,-2487.7,-2476.0,-16613.,-142.94,-20077.,-6375.8,-4361.8,-2797.9,66.782,2379.1,2169.3,1263.8,328.48,2603.2,1686.6,0.0000,6380.2,4449.7,4254.2,3660.4,0.0000,-380.25,-118.66,-77.574,-44.523,-83.181,-587.69,0.0000,-1069.5,-1585.9,-755.35,-1277.5
762.0000000000,94.936,2005.3,2069.8,1206.0,298.82,2405.4,972.09,1.5103,5273.1,2665.7,3354.0,1975.1,0.0000,-7218.0,-7140.9,-1462.5,-2486.6,-2471.6,-16610.,-142.81,-20074.,-6375.4,-4361.1,-2796.9,68.976,2390.8,2185.7,1267.2,335.09,2610.3,1686.6,2.0883,6383.8,4453.5,4259.6,3664.3,0.0000,-381.23,-119.18,-77.704,-44.678,-83.167,-587.69,-0.95605E-01,-1069.5,-1585.8,-755.36,-1277.4
763.0000000000,94.984,2006.7,2070.7,1204.1,298.94,2401.6,972.09,1.5262,5270.4,2665.8,3354.0,1975.3,0.0000,-7215.5,-7139.8,-1460.8,-2485.5,-2467.2,-16607.,-142.68,-20072.,-6374.9,-4360.3,-2796.0,66.877,2382.5,2172.4,1261.8,328.58,2597.1,1686.6,0.0000,6376.5,4449.7,4252.8,3658.0,0.0000,-380.71,-118.78,-77.556,-44.585,-82.827,-587.69,0.0000,-1069.3,-1585.6,-755.31,-1277.0
764.0000000000,94.944,2006.1,2070.3,1202.5,298.83,2397.5,972.09,1.5316,5267.3,2666.0,3354.1,1975.5,0.0000,-7213.0,-7138.8,-1459.1,-2484.4,-2462.9,-16604.,-142.55,-20069.,-6374.5,-4359.5,-2795.0,66.804,2379.9,2170.0,1259.0,328.19,2590.6,1686.6,0.0000,6372.5,4449.7,4252.8,3658.0,0.0000,-380.24,-118.62,-77.421,-44.536,-82.535,-587.69,0.0000,-1069.2,-1585.5,-755.29,-1276.8
765.0000000000,94.926,2004.5,2068.7,1200.7,298.74,2392.9,972.09,1.5321,5264.1,2666.1,3354.1,1975.7,0.0000,-7210.4,-7137.7,-1457.4,-2483.3,-2458.6,-16601.,-142.42,-20067.,-6374.0,-4358.8,-2794.1,66.730,2377.2,2167.6,1256.1,327.80,2584.0,1686.6,0.0000,6368.5,4449.7,4252.8,3658.0,0.0000,-379.78,-118.47,-77.285,-44.486,-82.243,-587.69,0.0000,-1069.1,-1585.3,-755.27,-1276.6
766.0000000000,94.878,2002.4,2066.9,1198.6,298.38,2387.5,972.02,1.5326,5260.8,2666.3,3354.1,1975.9,0.0000,-7207.7,-7136.5,-1455.6,-2482.2,-2454.3,-16599.,-142.29,-20064.,-6373.6,-4358.0,-2793.1,66.628,2373.6,2164.3,1252.9,327.28,2576.7,1686.6,0.0000,6364.2,4449.7,4252.8,3658.0,0.0000,-379.15,-118.26,-77.122,-44.418,-81.929,-587.69,0.0000,-1069.0,-1585.2,-755.26,-1276.4
767.0000000000,94.802,2000.1,2064.8,1196.3,297.96,2381.8,972.01,1.5330,5257.3,2666.5,3354.1,1976.1,0.0000,-7204.9,-7135.3,-1453.9,-2481.1,-2450.0,-16596.,-142.16,-20061.,-6373.1,-4357.3,-2792.2,66.545,2370.6,2161.6,1250.0,326.85,2570.1,1686.6,0.0000,6360.2,4449.7,4252.8,3658.0,0.0000,-378.63,-118.08,-76.980,-44.363,-81.636,-587.69,0.0000,-1068.9,-1585.0,-755.24,-1276.2
768.0000000000,94.881,1997.7,2062.5,1193.8,297.58,2376.0,972.01,1.5335,5253.9,2666.6,3354.1,1976.3,0.0000,-7202.1,-7134.1,-1452.2,-2480.0,-2445.6,-16593.,-142.03,-20059.,-6372.7,-4356.5,-2791.2,66.443,2367.0,2158.3,1246.8,326.33,2563.0,1686.6,0.0000,6355.9,4449.7,4252.8,3658.0,0.0000,-378.01,-117.88,-76.820,-44.296,-81.329,-587.69,0.0000,-1068.8,-1584.9,-755.22,-1276.0
769.0000000000,94.778,1995.0,2060.1,1191.0,297.13,2370.2,972.01,1.5340,5250.6,2666.8,3354.2,1976.5,0.0000,-7199.1,-7132.8,-1450.4,-2478.8,-2441.2,-16590.,-141.90,-20056.,-6372.2,-4355.8,-2790.3,66.324,2362.8,2154.5,1243.4,325.73,2555.5,1686.6,0.0000,6351.3,4449.7,4252.8,3658.0,0.0000,-377.28,-117.64,-76.641,-44.216,-81.005,-587.69,0.0000,-1068.7,-1584.7,-755.20,-1275.8
770.0000000000,94.636,1992.0,2057.3,1188.2,296.63,2364.8,972.02,1.5345,5248.0,2666.9,3354.2,1976.7,0.0000,-7196.1,-7131.4,-1448.6,-2477.7,-2436.8,-16588.,-141.78,-20053.,-6371.8,-4355.0,-2789.4,66.184,2357.8,2149.9,1239.6,325.02,2547.2,1686.6,0.0000,6346.3,4449.7,4252.8,3658.0,0.0000,-376.44,-117.36,-76.440,-44.123,-80.660,-587.69,0.0000,-1068.6,-1584.6,-755.18,-1275.6
771.0000000000,94.067,1988.6,2053.8,1185.4,296.06,2359.5,972.02,1.5350,5245.1,2666.8,3354.2,1976.9,0.0000,-7192.8,-7130.0,-1446.8,-2476.5,-2432.4,-16585.,-141.65,-20051.,-6371.3,-4354.3,-2788.4,66.044,2352.8,2145.4,1235.9,324.31,2539.0,1686.6,0.0000,6341.4,4449.7,4252.8,3658.0,0.0000,-375.59,-117.08,-76.239,-44.029,-80.316,-587.69,0.0000,-1068.5,-1584.4,-755.17,-1275.4
772.0000000000,93.845,1984.9,2050.0,1182.3,295.45,2353.7,972.01,1.5372,5241.9,2666.9,3354.2,1977.1,0.0000,-7189.4,-7128.5,-1444.9,-2475.4,-2427.9,-16582.,-141.52,-20048.,-6370.9,-4353.5,-2787.5,65.901,2347.7,2140.7,1232.0,323.59,2530.8,1686.6,0.0000,6336.3,4449.7,4252.8,3658.0,0.0000,-374.72,-116.79,-76.034,-43.934,-79.969,-587.69,0.0000,-1068.4,-1584.3,-755.15,-1275.2
773.0000000000,93.817,1981.4,2046.1,1179.2,294.85,2347.5,972.01,1.5467,5238.5,2667.1,3354.2,1977.3,0.0000,-7185.9,-7127.0,-1443.1,-2474.2,-2423.5,-16579.,-141.39,-20046.,-6370.4,-4352.7,-2786.5,65.759,2342.6,2136.1,1228.3,322.87,2522.6,1686.6,0.0000,6331.4,4449.7,4252.8,3658.0,0.0000,-373.86,-116.50,-75.833,-43.839,-79.626,-587.69,0.0000,-1068.3,-1584.1,-755.13,-1275.0
774.0000000000,93.743,1977.6,2042.3,1176.0,294.26,2340.9,971.85,1.5472,5234.8,2667.3,3354.3,1977.5,0.0000,-7182.3,-7125.4,-1441.2,-2473.0,-2419.0,-16576.,-141.26,-20043.,-6370.0,-4352.0,-2785.6,65.648,2338.7,2132.5,1225.0,322.31,2515.3,1686.6,0.0000,6327.0,4449.7,4252.8,3658.0,0.0000,-373.17,-116.27,-75.664,-43.765,-79.314,-587.69,0.0000,-1068.2,-1584.0,-755.11,-1274.8
775.0000000000,93.611,1974.1,2038.8,1172.7,293.71,2334.1,971.83,1.5476,5231.0,2667.4,3354.2,1977.7,0.0000,-7178.5,-7123.7,-1439.3,-2471.8,-2414.5,-16574.,-141.13,-20040.,-6369.5,-4351.2,-2784.6,65.521,2334.2,2128.4,1221.5,321.67,2507.7,1686.6,0.0000,6322.4,4449.7,4252.8,3658.0,0.0000,-372.39,-116.01,-75.479,-43.681,-78.988,-587.69,0.0000,-1068.1,-1583.8,-755.09,-1274.6
776.0000000000,93.624,1970.6,2035.4,1169.4,293.14,2327.8,971.83,1.5481,5227.0,2667.6,3354.2,1977.9,0.0000,-7174.7,-7122.1,-1437.4,-2470.7,-2410.0,-16571.,-141.00,-20038.,-6369.1,-4350.5,-2783.7,65.389,2329.5,2124.1,1217.9,321.00,2499.8,1686.6,0.0000,6317.6,4449.7,4252.8,3658.0,0.0000,-371.58,-115.74,-75.288,-43.593,-78.657,-587.69,0.0000,-1068.0,-1583.7,-755.08,-1274.4
777.0000000000,93.260,1967.1,2031.7,1166.1,292.59,2321.6,971.82,1.5486,5223.0,2667.7,3354.2,1978.1,0.0000,-7170.9,-7120.4,-1435.5,-2469.5,-2405.5,-16568.,-140.88,-20035.,-6368.6,-4349.7,-2782.8,65.266,2325.1,2120.1,1214.5,320.37,2492.2,1686.6,0.0000,6313.0,4449.7,4252.8,3658.0,0.0000,-370.82,-115.48,-75.106,-43.511,-78.333,-587.69,0.0000,-1067.9,-1583.5,-755.06,-1274.2
778.0000000000,93.119,1963.9,2028.3,1163.0,292.09,2315.0,971.80,1.5491,5219.1,2667.9,3354.2,1978.3,0.0000,-7166.9,-7118.7,-1433.6,-2468.3,-2400.9,-16565.,-140.75,-20032.,-6368.2,-4349.0,-2781.8,65.203,2322.8,2118.0,1211.8,320.04,2486.1,1686.6,0.0000,6309.3,4449.7,4252.8,3658.0,0.0000,-370.40,-115.33,-74.983,-43.468,-78.057,-587.69,0.0000,-1067.8,-1583.4,-755.04,-1274.0
779.0000000000,93.019,1961.2,2025.3,1159.9,291.65,2308.7,971.81,1.5496,5215.1,2668.1,3354.2,1978.5,0.0000,-7163.0,-7117.0,-1431.7,-2467.1,-2396.4,-16563.,-140.62,-20030.,-6367.7,-4348.2,-2780.9,65.107,2319.4,2114.9,1208.8,319.55,2479.4,1686.6,0.0000,6305.3,4449.7,4252.8,3658.0,0.0000,-369.80,-115.13,-74.832,-43.405,-77.765,-587.69,0.0000,-1067.7,-1583.3,-755.02,-1273.8
780.0000000000,92.910,1958.3,2022.4,1156.9,291.12,2302.2,971.81,1.5501,5211.2,2668.1,3354.3,1978.7,0.0000,-7159.0,-7115.3,-1429.8,-2465.9,-2391.9,-16560.,-140.49,-20027.,-6367.3,-4347.5,-2779.9,64.993,2315.3,2111.2,1205.6,318.97,2472.3,1686.6,0.0000,6301.0,4449.7,4252.8,3658.0,0.0000,-369.09,-114.89,-74.663,-43.329,-77.457,-587.69,0.0000,-1067.5,-1583.1,-755.01,-1273.6
781.0000000000,92.799,1955.1,2019.5,1154.0,290.60,2295.7,971.79,1.5506,5207.1,2668.3,3354.3,1978.9,0.0000,-7155.0,-7113.6,-1427.8,-2464.7,-2387.4,-16557.,-140.37,-20024.,-6366.8,-4346.7,-2779.0,64.862,2310.7,2107.0,1202.1,318.31,2464.6,1686.6,0.0000,6296.3,4449.7,4252.8,3658.0,0.0000,-368.28,-114.62,-74.475,-43.241,-77.132,-587.69,0.0000,-1067.4,-1583.0,-754.99,-1273.4
782.0000000000,92.843,1951.4,2015.8,1151.0,290.03,2289.1,971.76,1.5511,5203.1,2668.5,3354.3,1979.1,0.0000,-7150.9,-7111.8,-1425.9,-2463.5,-2382.9,-16554.,-140.24,-20022.,-6366.4,-4346.0,-2778.0,64.706,2305.1,2101.9,1198.1,317.52,2456.2,1686.6,0.0000,6291.2,4449.7,4252.8,3658.0,0.0000,-367.33,-114.30,-74.260,-43.137,-76.782,-587.69,0.0000,-1067.3,-1582.8,-754.97,-1273.1
783.0000000000,92.701,1947.4,2011.7,1148.0,289.41,2282.3,971.76,1.5516,5199.1,2668.6,3354.3,1979.3,0.0000,-7146.7,-7110.0,-1424.0,-2462.3,-2378.3,-16552.,-140.11,-20019.,-6365.9,-4345.2,-2777.1,64.552,2299.6,2096.9,1194.2,316.75,2447.7,1686.6,0.0000,6286.1,4449.7,4252.8,3658.0,0.0000,-366.39,-113.99,-74.047,-43.034,-76.434,-587.69,0.0000,-1067.2,-1582.7,-754.95,-1272.9
784.0000000000,92.551,1943.4,2007.6,1144.7,288.79,2275.5,971.76,1.5520,5195.0,2668.7,3354.3,1979.5,0.0000,-7142.3,-7108.1,-1422.0,-2461.0,-2373.8,-16549.,-139.98,-20017.,-6365.5,-4344.5,-2776.2,64.447,2295.9,2093.5,1191.1,316.21,2440.8,1686.6,0.0000,6282.0,4449.7,4252.8,3658.0,0.0000,-365.73,-113.76,-73.886,-42.965,-76.134,-587.69,0.0000,-1067.1,-1582.5,-754.93,-1272.7
785.0000000000,92.420,1940.1,2004.2,1141.3,288.28,2268.7,971.76,1.5525,5190.9,2668.9,3354.3,1979.7,0.0000,-7138.0,-7106.2,-1420.1,-2459.8,-2369.2,-16546.,-139.86,-20014.,-6365.0,-4343.7,-2775.2,64.379,2293.5,2091.3,1188.6,315.86,2435.1,1686.6,0.0000,6278.5,4449.7,4252.8,3658.0,0.0000,-365.27,-113.60,-73.766,-42.919,-75.873,-587.69,0.0000,-1067.0,-1582.4,-754.92,-1272.5
786.0000000000,92.312,1937.5,2001.4,1138.2,287.85,2262.1,971.77,1.5530,5187.0,2669.0,3354.4,1979.9,0.0000,-7133.7,-7104.4,-1418.1,-2458.6,-2364.6,-16543.,-139.73,-20011.,-6364.6,-4342.9,-2774.3,64.300,2290.7,2088.7,1186.0,315.45,2429.1,1686.6,0.0000,6274.9,4449.7,4252.8,3658.0,0.0000,-364.76,-113.42,-73.635,-42.867,-75.602,-587.69,0.0000,-1066.9,-1582.2,-754.90,-1272.3
787.0000000000,92.211,1934.8,1998.5,1135.3,287.44,2255.9,971.77,1.5535,5183.2,2669.1,3354.4,1980.1,0.0000,-7129.4,-7102.6,-1416.1,-2457.4,-2360.1,-16541.,-139.60,-20009.,-6364.1,-4342.2,-2773.3,64.184,2286.5,2084.9,1182.7,314.86,2421.9,1686.6,0.0000,6270.5,4449.7,4252.8,3658.0,0.0000,-364.03,-113.17,-73.463,-42.789,-75.295,-587.69,0.0000,-1066.8,-1582.1,-754.88,-1272.1
788.0000000000,92.103,1931.8,1995.5,1132.5,287.01,2249.7,971.77,1.5539,5179.4,2669.3,3354.4,1980.3,0.0000,-7125.0,-7100.7,-1414.2,-2456.1,-2355.5,-16538.,-139.48,-20006.,-6363.7,-4341.4,-2772.4,64.091,2283.2,2081.9,1179.8,314.39,2415.5,1686.6,0.0000,6266.6,4449.7,4252.8,3658.0,0.0000,-363.44,-112.96,-73.317,-42.727,-75.011,-587.69,0.0000,-1066.7,-1581.9,-754.86,-1271.9
789.0000000000,92.008,1929.4,1992.9,1129.6,286.68,2243.6,971.77,1.5544,5175.6,2669.4,3354.4,1980.5,0.0000,-7120.7,-7098.9,-1412.2,-2454.9,-2351.0,-16535.,-139.35,-20003.,-6363.2,-4340.7,-2771.5,64.095,2283.3,2082.0,1178.6,314.38,2412.4,1686.6,0.0000,6264.7,4449.7,4252.8,3658.0,0.0000,-363.39,-112.93,-73.278,-42.730,-74.834,-587.69,0.0000,-1066.6,-1581.8,-754.84,-1271.7
790.0000000000,91.958,1927.8,1990.9,1127.0,286.44,2237.7,971.77,1.5549,5171.9,2669.6,3354.4,1980.7,0.0000,-7116.4,-7097.1,-1410.3,-2453.7,-2346.4,-16532.,-139.23,-20000.,-6362.8,-4339.9,-2770.5,64.034,2281.2,2080.0,1176.3,314.06,2406.9,1686.6,0.0000,6261.4,4449.7,4252.8,3658.0,0.0000,-362.98,-112.78,-73.165,-42.689,-74.582,-587.69,0.0000,-1066.6,-1581.6,-754.83,-1271.5
791.0000000000,91.885,1926.0,1989.0,1124.6,286.14,2232.0,971.75,1.5554,5168.0,2669.7,3354.4,1980.9,0.0000,-7112.2,-7095.4,-1408.4,-2452.5,-2341.9,-16530.,-139.10,-19998.,-6362.3,-4339.2,-2769.6,63.943,2277.9,2077.1,1173.5,313.60,2400.7,1686.6,0.0000,6257.6,4449.7,4252.8,3658.0,0.0000,-362.39,-112.58,-73.023,-42.629,-74.305,-587.69,0.0000,-1066.5,-1581.5,-754.81,-1271.3
792.0000000000,91.806,1923.5,1986.5,1122.2,285.83,2226.3,971.73,1.5558,5164.3,2669.9,3354.4,1981.1,0.0000,-7108.0,-7093.6,-1406.5,-2451.3,-2337.4,-16527.,-138.98,-19995.,-6361.9,-4338.4,-2768.6,63.836,2274.1,2073.6,1170.4,313.06,2393.8,1686.6,0.0000,6253.5,4449.7,4252.8,3658.0,0.0000,-361.72,-112.35,-72.862,-42.558,-74.010,-587.69,0.0000,-1066.4,-1581.4,-754.79,-1271.1
793.0000000000,91.722,1920.6,1983.7,1119.6,285.41,2220.8,971.72,1.5500,5160.7,2670.0,3354.5,1981.3,0.0000,-7103.7,-7091.9,-1404.5,-2450.1,-2332.9,-16524.,-138.85,-19992.,-6361.4,-4337.7,-2767.7,63.704,2269.4,2069.3,1166.9,312.39,2386.3,1686.6,0.0000,6249.0,4449.7,4252.8,3658.0,0.0000,-360.91,-112.07,-72.676,-42.469,-73.694,-587.69,0.0000,-1066.3,-1581.2,-754.77,-1270.9
794.0000000000,91.607,1918.7,1981.6,1117.1,285.14,2215.4,971.69,1.5505,5157.1,2670.1,3354.5,1981.5,0.0000,-7099.4,-7090.1,-1402.6,-2448.9,-2328.4,-16521.,-138.73,-19990.,-6361.0,-4336.9,-2766.8,64.029,2276.2,2075.4,1168.6,313.40,2388.3,1686.6,0.18878,6250.3,4449.9,4253.0,3658.2,0.0000,-361.86,-112.36,-72.818,-42.590,-73.674,-587.69,-0.86410E-02,-1066.2,-1581.1,-754.75,-1270.7
795.0000000000,91.575,1919.0,1981.3,1114.7,285.21,2210.4,971.69,1.5509,5153.8,2670.3,3354.5,1981.7,0.0000,-7095.4,-7088.5,-1400.7,-2447.7,-2323.8,-16519.,-138.61,-19987.,-6360.5,-4336.2,-2765.8,63.811,2273.2,2072.8,1165.8,312.86,2382.2,1686.6,0.0000,6246.4,4449.7,4252.8,3658.0,0.0000,-361.38,-112.18,-72.692,-42.541,-73.408,-587.69,0.0000,-1066.1,-1580.9,-754.74,-1270.5
796.0000000000,91.303,1918.0,1980.4,1112.9,284.92,2205.6,971.69,1.5514,5150.5,2670.4,3354.5,1981.9,0.0000,-7091.4,-7086.9,-1398.9,-2446.5,-2319.4,-16516.,-138.48,-19984.,-6360.1,-4335.4,-2764.9,63.718,2269.9,2069.8,1162.9,312.38,2375.7,1686.6,0.0000,6242.5,4449.7,4252.8,3658.0,0.0000,-360.79,-111.98,-72.544,-42.478,-73.125,-587.69,0.0000,-1066.0,-1580.8,-754.72,-1270.3
797.0000000000,91.241,1916.3,1978.6,1111.0,284.83,2200.7,971.69,1.5518,5147.4,2670.6,3354.5,1982.1,0.0000,-7087.3,-7085.3,-1397.0,-2445.4,-2314.9,-16513.,-138.36,-19982.,-6359.6,-4334.7,-2764.0,63.692,2269.0,2068.9,1161.2,312.24,2371.6,1686.6,0.0000,6240.0,4449.7,4252.8,3658.0,0.0000,-360.58,-111.90,-72.474,-42.461,-72.920,-587.69,0.0000,-1065.9,-1580.6,-754.70,-1270.1
798.0000000000,91.229,1914.7,1976.7,1108.9,284.59,2195.7,971.66,1.5523,5144.3,2670.7,3354.5,1982.3,0.0000,-7083.3,-7083.7,-1395.1,-2444.2,-2310.5,-16510.,-138.23,-19979.,-6359.2,-4333.9,-2763.0,63.585,2265.2,2065.5,1158.1,311.69,2364.8,1686.6,0.0000,6235.9,4449.7,4252.8,3658.0,0.0000,-359.90,-111.67,-72.314,-42.390,-72.629,-587.69,0.0000,-1065.8,-1580.5,-754.68,-1269.9
799.0000000000,91.136,1912.5,1974.5,1106.8,284.17,2190.8,971.66,1.5553,5141.2,2670.8,3354.6,1982.5,0.0000,-7079.3,-7082.1,-1393.2,-2443.0,-2306.0,-16508.,-138.11,-19976.,-6358.7,-4333.2,-2762.1,63.491,2261.8,2062.4,1155.3,311.21,2358.6,1686.6,0.0000,6232.2,4449.7,4252.8,3658.0,0.0000,-359.31,-111.47,-72.169,-42.327,-72.355,-587.69,0.0000,-1065.7,-1580.4,-754.66,-1269.7
800.0000000000,91.044,1909.9,1971.4,1104.5,283.71,2185.6,971.62,1.5580,5138.1,2671.0,3354.6,1982.7,0.0000,-7075.1,-7080.4,-1391.3,-2441.8,-2301.5,-16505.,-137.99,-19974.,-6358.3,-4332.4,-2761.2,63.350,2256.8,2057.8,1151.7,310.50,2350.8,1686.6,0.0000,6227.5,4449.7,4252.8,3658.0,0.0000,-358.45,-111.18,-71.974,-42.233,-72.033,-587.69,0.0000,-1065.6,-1580.2,-754.65,-1269.5
801.0000000000,90.930,1906.6,1967.9,1102.0,283.17,2180.0,971.62,1.5584,5134.9,2671.1,3354.6,1982.9,0.0000,-7070.9,-7078.7,-1389.5,-2440.6,-2297.1,-16502.,-137.87,-19971.,-6357.8,-4331.7,-2760.2,63.211,2251.9,2053.3,1148.1,309.80,2343.1,1686.6,0.0000,6222.8,4449.7,4252.8,3658.0,0.0000,-357.59,-110.89,-71.780,-42.141,-71.713,-587.69,0.0000,-1065.5,-1580.1,-754.63,-1269.3
802.0000000000,90.797,1903.1,1964.5,1099.3,282.61,2174.1,971.58,1.5589,5131.6,2671.2,3354.6,1983.1,0.0000,-7066.6,-7077.0,-1387.6,-2439.4,-2292.6,-16499.,-137.74,-19968.,-6357.4,-4330.9,-2759.3,63.070,2246.8,2048.7,1144.5,309.10,2335.4,1686.6,0.0000,6218.1,4449.7,4252.8,3658.0,0.0000,-356.73,-110.61,-71.584,-42.047,-71.392,-587.69,0.0000,-1065.4,-1579.9,-754.61,-1269.1
803.0000000000,90.658,1899.4,1960.7,1096.4,281.91,2168.2,971.57,1.5593,5128.6,2671.3,3354.6,1983.3,0.0000,-7062.2,-7075.2,-1385.6,-2438.2,-2288.1,-16497.,-137.62,-19966.,-6356.9,-4330.1,-2758.4,62.923,2241.6,2044.0,1140.9,308.36,2327.5,1686.6,0.0000,6213.3,4449.7,4252.8,3658.0,0.0000,-355.83,-110.31,-71.383,-41.949,-71.067,-587.69,0.0000,-1065.3,-1579.8,-754.59,-1268.9
804.0000000000,90.508,1895.3,1956.7,1093.5,281.26,2162.4,971.56,1.5597,5125.4,2671.5,3354.6,1983.5,0.0000,-7057.7,-7073.4,-1383.7,-2436.9,-2283.6,-16494.,-137.50,-19963.,-6356.5,-4329.4,-2757.4,62.774,2236.3,2039.1,1137.2,307.61,2319.5,1686.6,0.0000,6208.5,4449.7,4252.8,3658.0,0.0000,-354.91,-110.00,-71.179,-41.849,-70.740,-587.69,0.0000,-1065.2,-1579.7,-754.57,-1268.8
805.0000000000,90.356,1891.4,1952.6,1090.3,280.62,2156.5,971.56,1.5602,5122.1,2671.6,3354.7,1983.7,0.0000,-7053.0,-7071.5,-1381.7,-2435.7,-2279.0,-16491.,-137.37,-19960.,-6356.0,-4328.6,-2756.5,62.627,2231.1,2034.4,1133.5,306.87,2311.6,1686.6,0.0000,6203.8,4449.7,4252.8,3658.0,0.0000,-354.01,-109.70,-70.978,-41.752,-70.417,-587.69,0.0000,-1065.1,-1579.5,-754.55,-1268.6
806.0000000000,90.304,1887.4,1948.5,1087.1,279.96,2150.3,971.56,1.5606,5118.6,2671.7,3354.7,1983.9,0.0000,-7048.3,-7069.6,-1379.8,-2434.4,-2274.5,-16489.,-137.25,-19958.,-6355.6,-4327.9,-2755.5,62.472,2225.5,2029.3,1129.7,306.09,2303.5,1686.6,0.0000,6198.9,4449.7,4252.8,3658.0,0.0000,-353.06,-109.38,-70.768,-41.648,-70.086,-587.69,0.0000,-1065.0,-1579.4,-754.54,-1268.4
807.0000000000,90.238,1883.5,1944.5,1083.9,279.25,2144.0,971.56,1.5610,5115.1,2671.9,3354.7,1984.1,0.0000,-7043.5,-7067.6,-1377.8,-2433.2,-2270.0,-16486.,-137.13,-19955.,-6355.1,-4327.1,-2754.6,62.387,2222.5,2026.6,1126.6,305.65,2296.5,1686.6,0.0000,6194.6,4449.7,4252.8,3658.0,0.0000,-352.51,-109.19,-70.619,-41.591,-69.787,-587.69,0.0000,-1064.9,-1579.3,-754.52,-1268.2
808.0000000000,90.115,1880.1,1940.7,1080.7,278.71,2138.4,971.56,1.5641,5111.4,2672.0,3354.7,1984.3,0.0000,-7038.7,-7065.7,-1375.8,-2432.0,-2265.4,-16483.,-137.01,-19952.,-6354.7,-4326.4,-2753.7,62.230,2216.9,2021.4,1122.7,304.86,2288.1,1686.6,0.0000,6189.5,4449.7,4252.8,3658.0,0.0000,-351.55,-108.87,-70.405,-41.486,-69.449,-587.69,0.0000,-1064.8,-1579.1,-754.50,-1268.0
809.0000000000,89.965,1877.3,1937.9,1077.5,278.26,2132.1,971.56,1.5837,5107.6,2672.1,3354.7,1984.5,0.0000,-7033.9,-7063.8,-1373.8,-2430.7,-2260.9,-16480.,-136.88,-19950.,-6354.2,-4325.6,-2752.7,62.502,2221.3,2025.5,1123.7,305.67,2289.0,1686.6,0.41481,6190.3,4450.1,4253.1,3658.3,0.0000,-352.14,-109.04,-70.492,-41.566,-69.395,-587.69,-0.18985E-01,-1064.7,-1579.0,-754.48,-1267.8
810.0000000000,89.954,1884.9,1944.2,1074.9,279.63,2127.2,971.57,1.6181,5103.9,2672.3,3354.7,1984.7,0.0000,-7030.0,-7062.3,-1371.9,-2429.6,-2256.5,-16478.,-136.77,-19947.,-6353.8,-4324.9,-2751.8,69.270,2290.8,2091.4,1147.0,316.99,2327.3,1686.6,11.027,6214.2,4453.7,4256.4,3661.7,0.0000,-362.12,-112.29,-72.144,-42.767,-70.457,-587.69,-0.50468,-1064.9,-1578.9,-754.48,-1267.7
811.0000000000,90.860,1911.0,1966.3,1074.7,283.76,2126.1,971.57,1.6245,5101.1,2672.4,3354.7,1984.9,0.0000,-7028.2,-7062.1,-1370.3,-2428.7,-2252.1,-16475.,-136.65,-19944.,-6353.3,-4324.1,-2750.9,221.93,2517.1,2330.3,1174.7,338.15,2363.5,1686.6,300.09,6241.8,4470.2,4272.3,3677.7,0.0000,-369.50,-118.70,-73.269,-43.700,-71.140,-587.69,-13.734,-1065.1,-1578.7,-754.55,-1268.1
812.0000000000,91.772,1939.0,1993.2,1078.8,287.49,2128.6,971.57,1.6282,5099.3,2672.5,3354.7,1985.1,0.0000,-7028.2,-7062.9,-1368.8,-2427.9,-2248.0,-16472.,-136.54,-19942.,-6352.9,-4323.4,-2750.0,66.142,2356.3,2148.5,1164.0,325.07,2348.6,1686.6,0.0000,6227.2,4453.4,4255.0,3660.1,0.0000,-373.45,-115.63,-73.771,-44.104,-70.979,-587.69,0.0000,-1064.8,-1578.6,-754.44,-1267.3
813.0000000000,92.628,1958.9,2013.0,1084.4,291.26,2131.8,971.56,1.6287,5098.2,2672.7,3354.8,1985.3,0.0000,-7029.2,-7064.1,-1367.5,-2427.3,-2244.2,-16469.,-136.42,-19939.,-6352.4,-4322.6,-2749.1,66.250,2360.1,2152.0,1160.8,324.24,2341.3,1686.6,0.0000,6221.3,4450.2,4253.1,3658.2,0.0000,-374.05,-115.82,-73.765,-44.168,-70.712,-587.69,0.0000,-1064.7,-1578.5,-754.41,-1267.0
814.0000000000,93.326,1968.2,2023.8,1088.4,293.18,2132.8,971.53,1.6292,5096.9,2672.8,3354.8,1985.4,0.0000,-7030.3,-7065.2,-1366.1,-2426.6,-2240.5,-16467.,-136.30,-19937.,-6352.0,-4321.9,-2748.1,66.206,2358.6,2150.6,1157.9,323.76,2334.5,1686.6,0.0000,6217.0,4449.8,4252.8,3658.0,0.0000,-373.79,-115.75,-73.648,-44.138,-70.433,-587.69,0.0000,-1064.6,-1578.3,-754.39,-1266.8
815.0000000000,93.656,1971.9,2028.7,1090.9,293.93,2131.8,971.49,1.6296,5095.0,2672.9,3354.8,1985.7,0.0000,-7031.0,-7066.0,-1364.8,-2425.8,-2236.7,-16464.,-136.18,-19934.,-6351.5,-4321.1,-2747.2,66.151,2356.6,2148.8,1155.8,323.43,2329.8,1686.6,0.0000,6214.1,4449.7,4252.8,3658.0,0.0000,-373.47,-115.66,-73.551,-44.100,-70.217,-587.69,0.0000,-1064.5,-1578.2,-754.37,-1266.7
816.0000000000,93.598,1973.2,2030.4,1092.0,293.86,2129.5,971.49,1.6301,5093.0,2673.1,3354.7,1985.8,0.0000,-7031.3,-7066.6,-1363.4,-2425.0,-2232.9,-16461.,-136.06,-19931.,-6351.1,-4320.4,-2746.3,66.053,2353.1,2145.6,1153.2,322.94,2324.2,1686.6,0.0000,6210.7,4449.7,4252.8,3658.0,0.0000,-372.91,-115.49,-73.412,-44.035,-69.973,-587.69,0.0000,-1064.4,-1578.1,-754.36,-1266.5
817.0000000000,93.538,1972.5,2031.2,1091.9,293.47,2126.5,971.49,1.6305,5091.7,2673.2,3354.7,1986.0,0.0000,-7031.2,-7066.9,-1362.1,-2424.1,-2229.0,-16459.,-135.94,-19929.,-6350.6,-4319.6,-2745.3,65.907,2347.9,2140.9,1150.1,322.21,2317.8,1686.6,0.0000,6206.9,4449.7,4252.8,3658.0,0.0000,-372.08,-115.24,-73.232,-43.938,-69.704,-587.69,0.0000,-1064.3,-1577.9,-754.34,-1266.3
818.0000000000,93.424,1970.9,2031.4,1091.1,292.93,2122.6,971.47,1.6310,5090.9,2673.3,3354.7,1986.2,0.0000,-7030.9,-7067.0,-1360.7,-2423.2,-2225.1,-16456.,-135.82,-19926.,-6350.2,-4318.9,-2744.4,65.724,2341.4,2135.0,1146.6,321.31,2310.7,1686.6,0.0000,6202.5,4449.7,4252.8,3658.0,0.0000,-371.03,-114.91,-73.016,-43.816,-69.413,-587.69,0.0000,-1064.2,-1577.8,-754.32,-1266.1
819.0000000000,93.585,1968.7,2029.8,1089.6,292.24,2119.6,971.46,1.6314,5091.9,2673.5,3354.7,1986.4,0.0000,-7030.3,-7066.8,-1359.2,-2422.2,-2221.1,-16453.,-135.70,-19923.,-6349.7,-4318.1,-2743.5,65.520,2334.1,2128.3,1142.8,320.31,2303.2,1686.6,0.0000,6198.0,4449.7,4252.8,3658.0,0.0000,-369.87,-114.55,-72.783,-43.680,-69.111,-587.69,0.0000,-1064.1,-1577.7,-754.30,-1265.9
820.0000000000,93.445,1964.9,2025.9,1088.0,291.44,2118.5,971.46,1.6318,5093.9,2673.6,3354.7,1986.6,0.0000,-7029.3,-7066.4,-1357.6,-2421.3,-2217.2,-16451.,-135.58,-19921.,-6349.3,-4317.4,-2742.6,65.308,2326.6,2121.5,1138.9,319.27,2295.6,1686.6,0.0000,6193.4,4449.7,4252.8,3658.0,0.0000,-368.65,-114.17,-72.542,-43.539,-68.805,-587.69,0.0000,-1064.0,-1577.5,-754.28,-1265.7
821.0000000000,93.375,1960.9,2020.9,1085.9,290.58,2117.7,971.46,1.6323,5094.8,2673.7,3354.8,1986.8,0.0000,-7027.7,-7065.9,-1355.9,-2420.2,-2213.2,-16448.,-135.46,-19918.,-6348.8,-4316.6,-2741.6,65.095,2319.0,2114.5,1135.1,318.23,2288.0,1686.6,0.0000,6188.9,4449.7,4252.8,3658.0,0.0000,-367.42,-113.79,-72.301,-43.397,-68.501,-587.69,0.0000,-1063.9,-1577.4,-754.27,-1265.5
822.0000000000,93.220,1956.9,2016.4,1083.3,289.68,2116.0,971.46,1.6327,5094.2,2673.9,3354.8,1987.0,0.0000,-7025.8,-7065.1,-1354.3,-2419.2,-2209.3,-16445.,-135.34,-19916.,-6348.4,-4315.9,-2740.7,64.873,2311.1,2107.3,1131.1,317.14,2280.1,1686.6,0.0000,6184.2,4449.7,4252.8,3658.0,0.0000,-366.14,-113.38,-72.051,-43.249,-68.190,-587.69,0.0000,-1063.8,-1577.3,-754.25,-1265.4
823.0000000000,92.997,1951.9,2011.5,1080.7,288.76,2111.9,971.46,1.6332,5092.3,2674.0,3354.8,1987.1,0.0000,-7023.4,-7064.3,-1352.6,-2418.2,-2205.3,-16442.,-135.23,-19913.,-6347.9,-4315.1,-2739.8,64.637,2302.7,2099.6,1126.9,315.99,2271.9,1686.6,0.0000,6179.2,4449.7,4252.8,3658.0,0.0000,-364.77,-112.95,-71.786,-43.091,-67.866,-587.69,0.0000,-1063.7,-1577.1,-754.23,-1265.2
824.0000000000,92.765,1946.5,2006.2,1077.8,287.83,2106.4,971.45,1.6336,5089.9,2674.1,3354.8,1987.3,0.0000,-7020.7,-7063.3,-1350.9,-2417.1,-2201.5,-16440.,-135.11,-19911.,-6347.5,-4314.4,-2738.8,64.432,2295.3,2093.0,1123.2,314.98,2264.5,1686.6,0.0000,6174.7,4449.7,4252.8,3658.0,0.0000,-363.57,-112.57,-71.552,-42.954,-67.568,-587.69,0.0000,-1063.6,-1577.0,-754.21,-1265.0
825.0000000000,92.545,1941.3,2001.8,1074.7,286.95,2100.3,971.45,1.6340,5086.8,2674.3,3354.8,1987.5,0.0000,-7017.8,-7062.2,-1349.1,-2416.0,-2197.6,-16437.,-134.99,-19908.,-6347.0,-4313.6,-2737.9,64.252,2289.0,2087.1,1119.8,314.10,2257.8,1686.6,0.0000,6170.7,4449.7,4252.8,3658.0,0.0000,-362.52,-112.23,-71.345,-42.835,-67.292,-587.69,0.0000,-1063.5,-1576.9,-754.19,-1264.8
826.0000000000,92.340,1936.5,1997.4,1071.2,286.14,2094.1,971.45,1.6345,5083.3,2674.4,3354.8,1987.7,0.0000,-7014.8,-7061.1,-1347.3,-2414.9,-2193.9,-16434.,-134.87,-19905.,-6346.6,-4312.9,-2737.0,64.107,2283.8,2082.4,1117.1,313.38,2252.3,1686.6,0.0000,6167.4,4449.7,4252.8,3658.0,0.0000,-361.66,-111.96,-71.176,-42.738,-67.052,-587.69,0.0000,-1063.4,-1576.7,-754.18,-1264.6
827.0000000000,92.339,1932.2,1992.5,1067.9,285.38,2088.3,971.45,1.6349,5079.6,2674.5,3354.9,1987.8,0.0000,-7011.6,-7059.8,-1345.5,-2413.8,-2190.2,-16432.,-134.75,-19903.,-6346.1,-4312.2,-2736.1,63.887,2276.0,2075.3,1113.1,312.31,2244.4,1686.6,0.0000,6162.6,4449.7,4252.8,3658.0,0.0000,-360.37,-111.55,-70.927,-42.592,-66.741,-587.69,0.0000,-1063.3,-1576.6,-754.16,-1264.4
828.0000000000,92.142,1926.8,1986.7,1064.6,284.52,2082.9,971.46,1.6353,5076.2,2674.7,3354.9,1988.0,0.0000,-7008.2,-7058.5,-1343.7,-2412.7,-2186.7,-16429.,-134.63,-19900.,-6345.7,-4311.4,-2735.1,63.661,2267.9,2067.9,1109.1,311.20,2236.6,1686.6,0.0000,6157.9,4449.7,4252.8,3658.0,0.0000,-359.04,-111.13,-70.674,-42.440,-66.431,-587.69,0.0000,-1063.2,-1576.5,-754.14,-1264.2
829.0000000000,92.119,1921.5,1981.1,1061.5,283.78,2077.3,971.46,1.6358,5072.9,2674.8,3354.9,1988.2,0.0000,-7004.6,-7057.0,-1341.9,-2411.6,-2183.3,-16426.,-134.52,-19898.,-6345.2,-4310.7,-2734.2,63.606,2265.9,2066.1,1107.4,310.92,2232.7,1686.6,0.0000,6155.6,4449.7,4252.8,3658.0,0.0000,-358.69,-111.01,-70.586,-42.404,-66.241,-587.69,0.0000,-1063.2,-1576.3,-754.12,-1264.1
830.0000000000,91.993,1917.1,1976.3,1058.8,283.15,2072.1,971.46,1.6362,5069.4,2675.1,3354.9,1988.4,0.0000,-7000.9,-7055.5,-1340.1,-2410.5,-2180.0,-16424.,-134.40,-19895.,-6344.8,-4309.9,-2733.3,63.370,2257.5,2058.5,1103.1,309.76,2224.3,1686.6,0.0000,6150.5,4449.7,4252.8,3658.0,0.0000,-357.30,-110.57,-70.319,-42.247,-65.914,-587.69,0.0000,-1063.1,-1576.2,-754.10,-1263.9
831.0000000000,91.728,1911.7,1970.8,1056.1,282.25,2066.4,971.46,1.6366,5065.5,2675.4,3354.9,1988.6,0.0000,-6996.9,-7053.9,-1338.2,-2409.3,-2176.9,-16421.,-134.29,-19892.,-6344.3,-4309.2,-2732.4,63.149,2249.6,2051.3,1099.0,308.68,2216.2,1686.6,0.0000,6145.6,4449.7,4252.8,3658.0,0.0000,-356.00,-110.16,-70.066,-42.099,-65.597,-587.69,0.0000,-1063.0,-1576.1,-754.08,-1263.7
832.0000000000,91.295,1906.4,1964.9,1053.3,281.54,2060.5,971.42,1.6370,5061.6,2675.5,3354.9,1988.7,0.0000,-6992.8,-7052.1,-1336.4,-2408.2,-2173.8,-16418.,-134.17,-19890.,-6343.9,-4308.4,-2731.4,63.010,2244.7,2046.8,1096.5,308.00,2211.2,1686.6,0.0000,6142.6,4449.7,4252.8,3658.0,0.0000,-355.16,-109.88,-69.907,-42.007,-65.374,-587.69,0.0000,-1062.9,-1575.9,-754.07,-1263.5
833.0000000000,91.140,1903.5,1962.1,1050.4,281.17,2054.5,971.42,1.6375,5058.0,2675.7,3354.9,1988.9,0.0000,-6988.8,-7050.5,-1334.6,-2407.0,-2170.9,-16416.,-134.06,-19887.,-6343.4,-4307.7,-2730.5,71.008,2265.4,2067.3,1105.3,313.04,2223.8,1686.6,15.428,6152.2,4455.0,4257.8,3662.9,0.0000,-356.91,-110.63,-70.225,-42.240,-65.567,-587.69,-0.70597,-1062.9,-1575.8,-754.07,-1263.5
834.0000000000,91.202,1904.6,1963.0,1048.2,281.37,2049.6,971.41,1.6379,5055.0,2675.7,3354.9,1989.1,0.0000,-6985.1,-7049.0,-1332.8,-2405.9,-2167.9,-16413.,-133.94,-19884.,-6343.0,-4306.9,-2729.6,63.245,2253.1,2054.4,1098.4,309.11,2213.4,1686.6,0.0000,6143.9,4449.7,4252.8,3658.0,0.0000,-356.37,-110.24,-70.092,-42.164,-65.282,-587.69,0.0000,-1062.8,-1575.7,-754.03,-1263.2
835.0000000000,91.140,1904.1,1963.6,1046.7,281.09,2045.5,971.40,1.6383,5051.8,2675.6,3355.0,1989.3,0.0000,-6981.5,-7047.5,-1331.1,-2404.8,-2164.9,-16410.,-133.83,-19882.,-6342.5,-4306.2,-2728.7,63.143,2249.4,2051.1,1095.5,308.59,2207.1,1686.6,0.0000,6140.1,4449.7,4252.8,3658.0,0.0000,-355.74,-110.03,-69.942,-42.095,-65.007,-587.69,0.0000,-1062.7,-1575.6,-754.01,-1263.0
836.0000000000,91.088,1902.6,1962.5,1045.2,281.20,2041.8,971.40,1.6487,5049.1,2675.8,3355.0,1989.5,0.0000,-6978.1,-7046.1,-1329.3,-2403.7,-2161.9,-16408.,-133.72,-19879.,-6342.1,-4305.4,-2727.8,63.205,2251.6,2053.1,1096.4,309.72,2212.7,1686.6,0.0000,6143.4,4451.2,4261.0,3665.9,0.0000,-356.03,-110.11,-69.984,-42.142,-64.956,-587.69,0.0000,-1062.6,-1575.4,-754.04,-1263.1
837.0000000000,91.148,1901.6,1961.3,1043.5,281.12,2037.6,971.39,1.6521,5046.2,2675.9,3355.0,1989.7,0.0000,-6974.7,-7044.6,-1327.6,-2402.6,-2158.9,-16405.,-133.61,-19877.,-6341.7,-4304.7,-2726.8,63.076,2247.0,2048.9,1093.0,308.24,2201.4,1686.6,0.0000,6136.6,4449.7,4252.8,3658.0,0.0000,-355.25,-109.86,-69.822,-42.051,-64.669,-587.69,0.0000,-1062.5,-1575.3,-753.98,-1262.6
838.0000000000,91.054,1902.0,1962.2,1042.5,281.13,2033.6,971.39,1.6525,5043.2,2676.0,3355.0,1989.8,0.0000,-6971.5,-7043.3,-1325.9,-2401.6,-2155.9,-16402.,-133.50,-19874.,-6341.2,-4303.9,-2725.9,86.595,2281.8,2077.0,1101.3,311.89,2206.1,1686.6,13.551,6143.8,4458.0,4261.9,3663.9,0.0000,-357.90,-110.93,-70.146,-42.376,-64.624,-587.69,-0.62008,-1062.5,-1575.2,-754.01,-1262.6
839.0000000000,91.265,1906.3,1966.4,1041.2,281.99,2030.1,971.39,1.6529,5040.5,2676.1,3355.0,1990.0,0.0000,-6968.7,-7042.2,-1324.2,-2400.5,-2152.9,-16400.,-133.39,-19871.,-6340.8,-4303.2,-2725.0,63.568,2264.6,2064.9,1092.6,310.49,2194.8,1686.6,0.0000,6132.5,4449.7,4252.8,3658.0,0.0000,-357.92,-110.67,-70.061,-42.379,-64.298,-587.69,0.0000,-1062.3,-1575.1,-753.94,-1262.3
840.0000000000,91.333,1908.2,1969.1,1040.1,281.99,2026.2,971.39,1.6534,5038.1,2676.2,3355.0,1990.2,0.0000,-6966.2,-7041.2,-1322.6,-2399.5,-2149.9,-16397.,-133.29,-19869.,-6340.3,-4302.5,-2724.1,63.490,2261.8,2062.4,1089.4,310.08,2187.2,1686.6,0.0000,6127.9,4449.7,4252.8,3658.0,0.0000,-357.43,-110.51,-69.910,-42.327,-63.986,-587.69,0.0000,-1062.2,-1574.9,-753.92,-1262.1
841.0000000000,91.334,1907.8,1968.8,1038.9,282.17,2021.6,971.39,1.6538,5035.9,2676.3,3355.1,1990.4,0.0000,-6963.6,-7040.1,-1321.0,-2398.5,-2146.8,-16394.,-133.18,-19866.,-6339.9,-4301.7,-2723.2,63.381,2257.9,2058.9,1086.1,309.52,2180.0,1686.6,0.0000,6123.6,4449.7,4252.8,3658.0,0.0000,-356.78,-110.30,-69.743,-42.254,-63.685,-587.69,0.0000,-1062.2,-1574.8,-753.90,-1261.9
842.0000000000,91.353,1905.5,1966.7,1036.9,281.88,2016.6,971.39,1.6542,5034.0,2676.4,3355.1,1990.5,0.0000,-6960.8,-7038.9,-1319.3,-2397.4,-2143.7,-16392.,-133.07,-19863.,-6339.4,-4301.0,-2722.2,63.231,2252.6,2054.0,1082.5,308.77,2172.4,1686.6,0.0000,6119.0,4449.7,4252.8,3658.0,0.0000,-355.89,-110.02,-69.543,-42.154,-63.372,-587.69,0.0000,-1062.1,-1574.7,-753.89,-1261.8
843.0000000000,91.183,1902.2,1963.5,1034.6,281.31,2012.1,971.36,1.6546,5032.0,2676.5,3355.1,1990.7,0.0000,-6957.8,-7037.7,-1317.6,-2396.4,-2140.6,-16389.,-132.97,-19861.,-6339.0,-4300.2,-2721.3,63.044,2245.9,2047.9,1078.6,307.84,2164.2,1686.6,0.0000,6114.0,4449.7,4252.8,3658.0,0.0000,-354.79,-109.67,-69.311,-42.029,-63.042,-587.69,0.0000,-1062.0,-1574.6,-753.87,-1261.6
844.0000000000,90.978,1899.0,1960.0,1032.0,280.77,2007.6,971.36,1.6551,5029.5,2676.6,3355.1,1990.9,0.0000,-6954.6,-7036.3,-1315.9,-2395.3,-2137.4,-16386.,-132.86,-19858.,-6338.5,-4299.5,-2720.4,63.046,2248.8,2048.3,1082.5,308.01,2168.4,1686.6,16.063,6121.3,4459.4,4261.6,3666.1,0.0000,-354.76,-109.66,-69.308,-42.032,-62.972,-587.69,-0.73499,-1062.0,-1574.4,-753.90,-1261.7
845.0000000000,90.903,1896.6,1957.5,1029.3,280.37,2003.5,971.36,1.6555,5027.4,2676.8,3355.1,1991.1,0.0000,-6951.4,-7034.9,-1314.2,-2394.2,-2134.3,-16384.,-132.76,-19855.,-6338.1,-4298.7,-2719.5,62.853,2239.1,2041.7,1074.7,306.90,2156.2,1686.6,0.0000,6109.2,4449.7,4252.8,3658.0,0.0000,-353.62,-109.29,-69.079,-41.902,-62.637,-587.69,0.0000,-1061.8,-1574.3,-753.83,-1261.2
846.0000000000,90.495,1892.9,1954.3,1026.9,279.64,1998.8,971.36,1.6559,5024.9,2676.9,3355.2,1991.2,0.0000,-6947.9,-7033.5,-1312.5,-2393.1,-2131.1,-16381.,-132.66,-19853.,-6337.6,-4298.0,-2718.6,62.644,2231.7,2034.9,1070.6,305.87,2148.1,1686.6,0.0000,6104.4,4449.7,4252.8,3658.0,0.0000,-352.40,-108.90,-68.834,-41.763,-62.311,-587.69,0.0000,-1061.7,-1574.2,-753.81,-1261.1
847.0000000000,90.282,1889.8,1950.8,1024.5,279.25,1994.4,971.36,1.6563,5022.3,2677.0,3355.2,1991.4,0.0000,-6944.4,-7032.0,-1310.8,-2392.0,-2127.9,-16378.,-132.55,-19850.,-6337.2,-4297.3,-2717.7,64.219,2251.4,2046.6,1085.2,310.70,2167.7,1686.6,46.212,6125.6,4471.7,4274.5,3678.1,0.0000,-353.15,-109.26,-69.002,-41.880,-62.473,-587.69,-2.1145,-1061.9,-1574.1,-753.91,-1261.5
848.0000000000,90.288,1888.8,1949.3,1022.2,279.12,1990.7,971.34,1.6567,5019.9,2677.2,3355.2,1991.6,0.0000,-6940.9,-7030.5,-1309.1,-2390.9,-2124.7,-16376.,-132.45,-19847.,-6336.7,-4296.5,-2716.7,62.664,2232.4,2035.6,1070.7,305.97,2148.0,1686.6,0.0000,6104.3,4449.7,4252.8,3658.0,0.0000,-352.41,-108.88,-68.846,-41.776,-62.144,-587.69,0.0000,-1061.6,-1573.9,-753.78,-1260.7
849.0000000000,90.177,1887.0,1947.3,1020.5,278.63,1986.8,971.32,1.6572,5017.0,2677.5,3355.2,1991.7,0.0000,-6937.4,-7029.1,-1307.4,-2389.8,-2121.6,-16373.,-132.35,-19845.,-6336.3,-4295.8,-2715.8,62.555,2228.5,2032.0,1068.0,305.42,2142.2,1686.6,0.0000,6100.8,4449.7,4252.8,3658.0,0.0000,-351.75,-108.66,-68.697,-41.703,-61.887,-587.69,0.0000,-1061.5,-1573.8,-753.76,-1260.6
850.0000000000,89.935,1884.4,1944.2,1018.9,278.37,1982.9,971.32,1.6576,5013.9,2677.7,3355.2,1991.9,0.0000,-6933.8,-7027.7,-1305.7,-2388.7,-2118.4,-16371.,-132.24,-19842.,-6335.8,-4295.0,-2714.9,62.404,2223.1,2027.1,1064.7,304.67,2135.5,1686.6,0.0000,6096.7,4449.7,4252.8,3658.0,0.0000,-350.85,-108.38,-68.509,-41.603,-61.604,-587.69,0.0000,-1061.4,-1573.7,-753.74,-1260.4
851.0000000000,89.713,1880.6,1940.7,1016.6,277.80,1978.4,971.32,1.6580,5010.9,2677.9,3355.2,1992.1,0.0000,-6930.1,-7026.2,-1304.1,-2387.6,-2115.2,-16368.,-132.14,-19839.,-6335.4,-4294.3,-2714.0,62.241,2217.3,2021.8,1061.3,303.86,2128.5,1686.6,0.0000,6092.5,4449.7,4252.8,3658.0,0.0000,-349.88,-108.06,-68.309,-41.494,-61.314,-587.69,0.0000,-1061.3,-1573.6,-753.72,-1260.2
852.0000000000,89.644,1876.5,1936.4,1014.5,277.15,1973.2,971.29,1.6584,5007.6,2677.9,3355.2,1992.3,0.0000,-6926.1,-7024.6,-1302.4,-2386.4,-2112.0,-16365.,-132.04,-19836.,-6334.9,-4293.6,-2713.1,62.056,2210.7,2015.8,1057.7,302.95,2121.1,1686.6,0.0000,6088.0,4449.7,4252.8,3658.0,0.0000,-348.78,-107.71,-68.088,-41.371,-61.009,-587.69,0.0000,-1061.2,-1573.4,-753.70,-1260.0
853.0000000000,89.582,1871.8,1931.8,1012.0,276.41,1967.9,971.21,1.6588,5004.4,2677.9,3355.3,1992.4,0.0000,-6922.1,-7023.5,-1300.7,-2385.3,-2108.7,-16363.,-131.93,-19834.,-6334.5,-4292.8,-2712.2,61.863,2203.8,2009.5,1053.9,302.00,2113.4,1686.6,0.0000,6083.4,4449.7,4252.8,3658.0,0.0000,-347.64,-107.35,-67.859,-41.242,-60.700,-587.69,0.0000,-1061.1,-1573.3,-753.69,-1259.9
854.0000000000,89.397,1866.6,1926.8,1009.3,275.62,1962.7,971.18,1.6592,5001.5,2678.0,3355.3,1992.6,0.0000,-6917.8,-7022.4,-1299.0,-2384.1,-2105.5,-16360.,-131.83,-19831.,-6334.0,-4292.1,-2711.3,61.656,2196.5,2002.8,1049.9,300.99,2105.5,1686.6,0.0000,6078.6,4449.7,4252.8,3658.0,0.0000,-346.42,-106.96,-67.618,-41.104,-60.382,-587.69,0.0000,-1061.0,-1573.2,-753.67,-1259.7
855.0000000000,89.198,1861.4,1921.3,1006.4,274.78,1957.1,971.19,1.6596,4998.5,2678.1,3355.3,1992.8,0.0000,-6913.4,-7021.1,-1297.3,-2382.9,-2102.2,-16357.,-131.72,-19828.,-6333.6,-4291.3,-2710.3,61.450,2189.1,1996.1,1046.1,299.97,2097.8,1686.6,0.0000,6074.0,4449.7,4252.8,3658.0,0.0000,-345.21,-106.57,-67.381,-40.967,-60.072,-587.69,0.0000,-1060.9,-1573.1,-753.65,-1259.5
856.0000000000,88.741,1856.0,1915.7,1003.2,273.92,1951.3,971.19,1.6668,4995.5,2678.3,3355.3,1992.9,0.0000,-6908.8,-7019.7,-1295.6,-2381.8,-2098.8,-16355.,-131.62,-19826.,-6333.1,-4290.6,-2709.4,61.245,2181.8,1989.5,1042.2,298.96,2089.9,1686.6,0.0000,6069.3,4449.7,4252.8,3658.0,0.0000,-343.99,-106.18,-67.141,-40.830,-59.755,-587.69,0.0000,-1060.8,-1572.9,-753.63,-1259.4
857.0000000000,88.518,1850.4,1910.0,1000.1,272.97,1945.8,971.19,1.6763,4993.0,2678.4,3355.3,1993.1,0.0000,-6904.0,-7018.0,-1293.9,-2380.6,-2095.5,-16352.,-131.52,-19823.,-6332.7,-4289.9,-2708.5,61.030,2174.2,1982.5,1038.2,297.91,2082.0,1686.6,0.0000,6064.5,4449.7,4252.8,3658.0,0.0000,-342.72,-105.77,-66.894,-40.687,-59.438,-587.69,0.0000,-1060.7,-1572.8,-753.61,-1259.2
858.0000000000,88.473,1845.0,1904.0,996.70,272.01,1940.4,971.19,1.6768,4990.1,2678.5,3355.4,1993.3,0.0000,-6899.1,-7016.2,-1292.2,-2379.3,-2092.1,-16349.,-131.42,-19820.,-6332.2,-4289.1,-2707.6,60.801,2166.0,1975.0,1033.9,296.79,2073.5,1686.6,0.0000,6059.4,4449.7,4252.8,3658.0,0.0000,-341.37,-105.34,-66.630,-40.534,-59.104,-587.69,0.0000,-1060.6,-1572.7,-753.60,-1259.0
859.0000000000,88.249,1839.0,1897.9,993.26,271.08,1934.7,971.19,1.6808,4986.9,2678.6,3355.4,1993.4,0.0000,-6894.0,-7014.2,-1290.5,-2378.1,-2088.7,-16347.,-131.32,-19818.,-6331.8,-4288.4,-2706.7,60.576,2158.0,1967.7,1029.7,295.68,2065.1,1686.6,0.0000,6054.3,4449.7,4252.8,3658.0,0.0000,-340.04,-104.91,-66.370,-40.384,-58.772,-587.69,0.0000,-1060.5,-1572.6,-753.58,-1258.9
860.0000000000,88.023,1832.8,1891.5,989.83,270.14,1928.4,971.19,1.6856,4983.4,2678.7,3355.4,1993.6,0.0000,-6888.7,-7012.1,-1288.8,-2376.9,-2085.3,-16344.,-131.21,-19815.,-6331.3,-4287.6,-2705.8,60.356,2150.2,1960.6,1025.6,294.60,2056.9,1686.6,0.0000,6049.3,4449.7,4252.8,3658.0,0.0000,-338.74,-104.49,-66.116,-40.237,-58.446,-587.69,0.0000,-1060.4,-1572.4,-753.56,-1258.7
861.0000000000,87.799,1839.3,1897.0,986.73,271.32,1923.3,971.18,1.6860,4979.9,2678.8,3355.4,1993.7,0.0000,-6884.4,-7010.5,-1287.2,-2375.7,-2081.9,-16341.,-131.12,-19812.,-6330.9,-4286.9,-2704.9,79.730,2290.2,2071.3,1070.9,311.54,2134.2,1686.6,40.744,6099.7,4459.2,4262.2,3667.1,0.0000,-353.72,-109.60,-68.803,-42.039,-60.456,-587.69,-1.8641,-1060.8,-1572.3,-753.59,-1258.8
862.0000000000,88.883,1877.3,1929.2,1000.3,277.67,1972.6,971.14,1.6864,4982.7,2679.0,3355.4,1993.9,0.0000,-6883.3,-7010.6,-1287.7,-2374.9,-2080.2,-16339.,-131.03,-19809.,-6330.4,-4286.2,-2704.0,446.46,3364.3,2568.5,1755.3,350.45,3837.3,1686.7,781.29,7136.9,4481.7,4292.9,3691.2,0.0000,-368.16,-122.58,-92.215,-43.669,-110.01,-587.69,-35.745,-1068.2,-1572.2,-753.73,-1259.4
863.0000000000,90.369,1925.8,1974.8,1103.3,283.89,2197.5,971.10,1.6869,5037.5,2679.1,3355.4,1994.1,0.0000,-6885.4,-7012.6,-1292.3,-2374.5,-2083.1,-16336.,-130.94,-19807.,-6330.0,-4285.4,-2703.1,412.27,2948.9,2387.4,2077.8,376.95,4547.3,1687.8,932.39,7581.3,4544.6,4354.1,3745.7,0.0000,-376.49,-120.42,-101.44,-44.844,-128.97,-587.71,-42.657,-1071.7,-1572.1,-754.04,-1261.0
864.0000000000,91.992,1968.0,2015.7,1303.0,303.25,2532.6,971.10,1.6873,5124.6,2679.2,3355.5,1994.3,0.0000,-6889.8,-7015.8,-1297.7,-2374.3,-2092.3,-16334.,-130.85,-19806.,-6329.5,-4284.7,-2702.2,68.043,2424.0,2210.3,2038.2,348.62,4467.8,1689.3,419.28,7547.4,4614.8,4415.7,3812.2,0.0000,-381.82,-117.84,-102.57,-45.377,-129.50,-587.73,-19.182,-1071.1,-1572.0,-754.34,-1262.9
865.0000000000,93.723,1998.4,2046.6,1463.8,311.98,2808.6,971.05,1.6878,5227.0,2679.4,3355.9,1994.4,0.0000,-6895.5,-7019.3,-1306.6,-2374.1,-2108.4,-16331.,-130.76,-19806.,-6329.1,-4284.0,-2701.3,68.361,2435.3,2220.6,1994.5,349.32,4474.1,1686.6,102.58,7526.4,4468.8,4267.1,3674.3,0.0000,-383.64,-118.43,-103.03,-45.584,-130.27,-587.69,-4.6930,-1070.7,-1571.8,-753.55,-1258.4
866.0000000000,94.745,2018.9,2069.4,1619.3,315.61,2981.9,971.02,1.6882,5304.9,2679.7,3355.8,1994.6,0.0000,-6901.4,-7022.7,-1317.1,-2373.8,-2121.0,-16328.,-130.67,-19805.,-6328.7,-4283.2,-2700.4,255.29,3058.0,2557.7,2195.4,436.82,4734.6,1695.2,372.86,7739.4,4629.1,4425.9,3827.3,0.0000,-388.66,-126.41,-104.93,-46.572,-134.62,-587.82,-17.058,-1073.3,-1571.7,-754.36,-1263.0
867.0000000000,95.699,2050.8,2100.5,1715.5,321.35,3125.1,970.99,1.6886,5363.8,2679.9,3356.5,1995.3,0.0000,-6908.6,-7026.8,-1328.9,-2373.7,-2131.1,-16326.,-130.58,-19804.,-6328.2,-4282.5,-2699.5,1263.0,3453.5,3307.0,2245.5,499.93,4787.7,1717.3,393.28,7782.4,4643.9,4442.9,3844.3,0.0000,-406.43,-145.66,-107.41,-48.916,-136.09,-588.17,-17.992,-1073.7,-1571.6,-754.43,-1263.4
868.0000000000,97.667,2103.3,2149.0,1795.2,329.05,3225.8,970.98,1.6891,5468.6,2679.8,3357.3,1998.2,0.0000,-6918.5,-7032.3,-1344.8,-2373.8,-2140.1,-16323.,-130.49,-19803.,-6327.8,-4281.8,-2698.6,73.412,2615.3,2384.7,2074.5,427.87,4613.1,1686.6,0.0000,7605.6,4458.6,4259.0,3662.8,0.0000,-412.24,-127.41,-108.26,-49.284,-135.58,-587.69,0.0000,-1071.2,-1571.5,-753.45,-1257.6
869.0000000000,98.889,2140.6,2190.0,1841.7,333.43,3309.4,970.98,4.1446,5607.6,2682.5,3358.8,1999.8,0.0000,-6929.7,-7038.4,-1357.0,-2374.0,-2147.9,-16321.,-130.41,-19803.,-6327.3,-4281.0,-2697.7,73.483,2617.8,2387.0,2063.4,376.63,4600.4,1686.6,0.0000,7594.6,4450.8,4253.3,3658.3,0.0000,-412.76,-127.64,-108.31,-49.014,-135.86,-587.69,0.0000,-1071.0,-1571.4,-753.40,-1257.3
870.0000000000,99.856,2158.6,2210.6,1859.5,337.02,3509.8,970.98,12.665,5839.2,2683.8,3360.6,1998.2,0.0000,-6940.6,-7043.8,-1367.1,-2374.1,-2154.7,-16319.,-130.32,-19803.,-6326.9,-4280.3,-2696.8,73.338,2612.6,2382.3,2060.3,372.21,4598.7,1686.6,0.0000,7592.3,4449.7,4252.8,3658.0,0.0000,-412.07,-127.48,-108.22,-48.894,-136.19,-587.69,0.0000,-1071.0,-1571.3,-753.38,-1257.1
871.0000000000,100.45,2171.2,2225.1,1865.8,338.86,3720.9,970.98,18.842,5996.8,2684.3,3360.4,1998.0,0.0000,-6951.1,-7048.8,-1375.6,-2374.1,-2160.8,-16316.,-130.23,-19803.,-6326.5,-4279.6,-2696.0,558.31,3103.6,2832.5,2251.6,536.81,4786.4,1686.6,0.0000,7694.1,4449.7,4252.8,3658.0,0.0000,-418.41,-138.19,-108.87,-50.527,-137.45,-587.69,0.0000,-1072.5,-1571.2,-753.36,-1256.9
872.0000000000,101.08,2190.0,2243.2,1880.4,340.88,3859.7,970.98,29.703,6094.3,2684.1,3358.9,1998.4,0.0000,-6961.4,-7053.8,-1382.9,-2374.1,-2166.4,-16314.,-130.14,-19803.,-6326.1,-4278.9,-2695.1,74.694,2660.9,2426.3,2066.6,378.25,4600.0,1686.6,0.0000,7592.8,4449.7,4252.8,3658.0,0.0000,-419.97,-130.03,-109.13,-49.796,-136.83,-587.69,0.0000,-1071.0,-1571.0,-753.35,-1256.8
873.0000000000,101.34,2204.7,2258.0,1905.3,341.87,3912.5,970.99,22.565,6145.7,2686.9,3358.1,1998.3,0.0000,-6971.3,-7058.7,-1389.6,-2374.0,-2171.7,-16312.,-130.05,-19804.,-6325.8,-4278.2,-2694.2,74.627,2658.6,2424.2,2066.6,377.93,4600.7,1686.6,0.0000,7593.3,4449.7,4252.8,3658.0,0.0000,-419.76,-130.01,-109.10,-49.752,-137.15,-587.69,0.0000,-1071.1,-1570.9,-753.33,-1256.6
874.0000000000,101.59,2212.5,2267.5,1922.6,342.86,3926.4,970.99,18.983,6172.5,2686.1,3358.7,1998.0,0.0000,-6980.6,-7063.2,-1395.6,-2374.0,-2176.9,-16310.,-129.96,-19805.,-6325.5,-4277.5,-2693.3,74.689,2769.5,2426.2,2202.4,378.23,4644.8,1686.6,204.58,7731.9,4593.5,4301.0,3712.8,0.0000,-420.43,-130.21,-109.15,-49.793,-137.67,-587.69,-9.3590,-1073.1,-1570.8,-753.57,-1258.2
875.0000000000,101.77,2218.1,2273.9,1924.8,343.02,3929.0,970.99,22.359,6173.9,2685.6,3358.0,1997.9,0.0000,-6989.4,-7067.2,-1401.1,-2373.8,-2181.9,-16308.,-129.88,-19806.,-6325.2,-4276.8,-2692.4,74.442,2651.9,2418.1,2066.4,377.08,4602.2,1686.6,0.0000,7594.2,4449.7,4252.8,3658.0,0.0000,-419.01,-129.86,-109.00,-49.628,-137.75,-587.69,0.0000,-1071.1,-1570.7,-753.30,-1256.3
876.0000000000,101.63,2217.4,2274.4,1926.8,342.38,3950.3,971.00,20.789,6176.0,2684.8,3357.5,1998.0,0.0000,-6997.2,-7070.9,-1406.2,-2373.6,-2186.9,-16306.,-129.79,-19807.,-6324.9,-4276.1,-2691.5,74.277,2646.1,2412.8,2065.9,376.32,4602.8,1686.6,0.0000,7594.6,4449.7,4252.8,3658.0,0.0000,-418.22,-129.65,-108.89,-49.518,-138.04,-587.69,0.0000,-1071.1,-1570.6,-753.29,-1256.2
877.0000000000,101.75,2215.9,2273.6,1927.4,341.60,3987.4,971.00,26.611,6203.1,2683.8,3357.5,1998.2,0.0000,-7004.1,-7074.0,-1411.0,-2373.3,-2192.5,-16304.,-129.70,-19807.,-6324.5,-4275.5,-2690.7,73.921,2633.4,2401.2,2064.5,374.65,4603.1,1686.6,0.0000,7594.9,4449.7,4252.8,3658.0,0.0000,-416.33,-129.10,-108.66,-49.280,-138.31,-587.69,0.0000,-1071.1,-1570.5,-753.27,-1256.0
878.0000000000,101.54,2212.7,2270.5,1933.5,340.35,4028.8,971.00,26.847,6222.9,2683.6,3357.3,1998.1,0.0000,-7010.0,-7076.7,-1415.4,-2373.0,-2198.2,-16302.,-129.61,-19808.,-6324.1,-4274.8,-2689.8,73.556,2620.4,2389.4,2063.1,372.96,4603.7,1686.6,0.0000,7595.3,4449.7,4252.8,3658.0,0.0000,-414.39,-128.52,-108.43,-49.037,-138.59,-587.69,0.0000,-1071.1,-1570.4,-753.26,-1255.9
879.0000000000,101.49,2217.3,2274.7,1943.4,341.05,4047.0,970.97,22.707,6223.2,2683.6,3357.1,1998.2,0.0000,-7015.8,-7079.4,-1419.6,-2372.6,-2203.9,-16301.,-129.52,-19809.,-6323.8,-4274.1,-2688.9,679.79,3510.0,3040.4,2245.3,506.45,4778.9,1686.6,748.41,7759.5,4594.9,4393.1,3785.9,0.0000,-425.80,-144.33,-109.78,-50.982,-140.07,-587.69,-34.236,-1073.5,-1570.3,-753.98,-1259.7
880.0000000000,102.21,2240.3,2293.4,1945.2,344.14,4060.7,970.96,18.212,6227.1,2683.9,3357.0,1998.4,0.0000,-7023.0,-7083.0,-1423.6,-2372.5,-2209.5,-16299.,-129.44,-19810.,-6323.4,-4273.4,-2688.0,75.836,2701.6,2463.4,2082.4,384.83,4624.5,1686.6,0.0000,7608.3,4452.7,4257.4,3662.1,0.0000,-427.49,-132.65,-110.17,-50.564,-139.64,-587.69,0.0000,-1071.3,-1570.2,-753.25,-1255.7
881.0000000000,102.81,2268.0,2322.3,1949.7,348.30,4063.8,970.97,16.968,6250.2,2684.1,3357.0,1998.4,0.0000,-7031.8,-7087.4,-1427.7,-2372.5,-2215.1,-16297.,-129.35,-19811.,-6323.0,-4272.7,-2687.1,1135.3,3487.5,3221.1,2277.5,545.34,4809.8,1686.6,477.77,7785.6,4616.2,4416.3,3814.8,0.0000,-442.41,-151.49,-111.92,-53.091,-141.08,-587.69,-21.855,-1073.8,-1570.0,-754.07,-1260.3
882.0000000000,104.69,2309.9,2358.9,1955.1,355.21,4073.8,970.97,22.277,6258.7,2684.3,3357.2,1998.6,0.0000,-7043.0,-7093.0,-1431.6,-2372.8,-2220.8,-16295.,-129.27,-19811.,-6322.6,-4272.1,-2686.2,79.248,2823.2,2574.3,2102.2,406.19,4637.0,1686.6,0.0000,7616.6,4451.1,4253.6,3659.5,0.0000,-447.08,-138.89,-112.63,-52.872,-140.55,-587.69,0.0000,-1071.3,-1569.9,-753.20,-1255.3
883.0000000000,105.69,2337.5,2387.0,1961.0,358.70,4094.5,970.97,18.933,6275.1,2684.4,3357.4,2000.0,0.0000,-7054.7,-7098.9,-1435.4,-2373.1,-2226.8,-16293.,-129.18,-19812.,-6322.2,-4271.4,-2685.3,79.271,2824.0,2575.0,2101.7,399.95,4639.2,1686.6,0.0000,7615.8,4449.7,4252.8,3658.1,0.0000,-447.40,-139.08,-112.68,-52.848,-140.87,-587.69,0.0000,-1071.3,-1569.8,-753.18,-1255.1
884.0000000000,106.65,2348.8,2398.4,1966.7,361.02,4098.2,970.97,16.317,6281.4,2684.4,3357.3,2000.6,0.0000,-7065.8,-7104.2,-1439.1,-2373.3,-2232.6,-16292.,-129.09,-19813.,-6321.8,-4270.7,-2684.5,79.076,2817.0,2568.7,2101.6,398.95,4641.3,1686.6,0.0000,7617.1,4449.7,4252.8,3658.0,0.0000,-446.49,-138.87,-112.58,-52.717,-141.18,-587.69,0.0000,-1071.4,-1569.7,-753.16,-1254.9
885.0000000000,106.95,2349.8,2404.5,1969.6,361.06,4119.6,970.98,18.919,6288.8,2686.5,3358.0,2000.5,0.0000,-7075.8,-7108.8,-1442.5,-2373.4,-2238.2,-16290.,-129.01,-19813.,-6321.4,-4270.0,-2683.6,78.790,2806.9,2559.4,2102.6,397.66,4647.1,1686.6,0.0000,7620.6,4449.7,4252.8,3658.0,0.0000,-445.06,-138.49,-112.47,-52.527,-141.60,-587.69,0.0000,-1071.4,-1569.6,-753.15,-1254.8
886.0000000000,107.52,2347.6,2406.0,1971.3,360.10,4138.1,970.98,26.370,6310.8,2688.0,3359.0,2000.2,0.0000,-7084.7,-7112.6,-1445.7,-2373.3,-2243.5,-16289.,-128.92,-19814.,-6321.0,-4269.4,-2682.7,78.458,2795.0,2548.6,2104.0,396.16,4654.5,1686.6,0.0000,7625.2,4449.7,4252.8,3658.0,0.0000,-443.35,-138.02,-112.34,-52.305,-142.07,-587.69,0.0000,-1071.4,-1569.5,-753.13,-1254.6
887.0000000000,107.02,2343.4,2404.4,1973.6,358.80,4142.3,970.97,31.036,6347.2,2689.7,3358.8,2000.5,0.0000,-7092.8,-7115.8,-1448.7,-2373.1,-2248.6,-16287.,-128.83,-19814.,-6320.6,-4268.7,-2681.8,78.098,2782.2,2536.9,2104.5,394.51,4660.0,1686.6,0.0000,7628.6,4449.7,4252.8,3658.0,0.0000,-441.47,-137.49,-112.18,-52.065,-142.46,-587.69,0.0000,-1071.5,-1569.4,-753.12,-1254.5
888.0000000000,106.68,2337.4,2400.0,1976.0,357.47,4155.0,970.97,28.463,6354.1,2689.2,3358.1,2001.0,0.0000,-7100.1,-7118.4,-1451.6,-2372.9,-2253.7,-16286.,-128.74,-19815.,-6320.3,-4268.0,-2680.9,77.725,2768.9,2524.8,2104.4,392.80,4664.0,1686.6,0.0000,7631.1,4449.7,4252.8,3658.0,0.0000,-439.51,-136.93,-111.98,-51.816,-142.78,-587.69,0.0000,-1071.5,-1569.3,-753.10,-1254.3
889.0000000000,106.28,2331.2,2393.6,1979.0,356.05,4173.8,970.98,23.216,6366.4,2689.1,3357.7,2000.9,0.0000,-7106.3,-7120.4,-1454.4,-2372.6,-2258.9,-16284.,-128.65,-19815.,-6320.0,-4267.4,-2680.1,77.341,2755.2,2512.3,2103.7,391.03,4666.5,1686.6,0.0000,7632.7,4449.7,4252.8,3658.0,0.0000,-437.46,-136.33,-111.76,-51.561,-143.06,-587.69,0.0000,-1071.5,-1569.2,-753.09,-1254.2
890.0000000000,105.31,2323.1,2388.7,1981.2,354.53,4190.2,970.98,25.203,6374.4,2687.7,3358.4,2000.7,0.0000,-7111.7,-7122.0,-1457.0,-2372.2,-2265.9,-16283.,-128.56,-19816.,-6319.6,-4266.8,-2679.2,76.954,2741.4,2499.7,2102.5,389.23,4667.5,1686.6,0.0000,7633.4,4449.7,4252.8,3658.0,0.0000,-435.39,-135.71,-111.52,-51.303,-143.28,-587.69,0.0000,-1071.6,-1569.0,-753.07,-1254.0
891.0000000000,104.93,2314.6,2380.8,1981.8,353.00,4195.2,970.98,27.221,6376.4,2688.0,3358.0,2001.2,0.0000,-7116.1,-7123.2,-1459.6,-2371.8,-2272.9,-16281.,-128.48,-19816.,-6319.3,-4266.1,-2678.3,76.562,2727.5,2487.0,2100.6,387.40,4667.2,1686.6,0.0000,7633.3,4449.7,4252.8,3658.0,0.0000,-433.27,-135.08,-111.26,-51.042,-143.46,-587.69,0.0000,-1071.6,-1568.9,-753.06,-1253.9
892.0000000000,104.53,2306.3,2372.4,1981.6,351.37,4209.1,970.98,28.454,6378.5,2688.3,3357.8,2001.2,0.0000,-7119.8,-7124.0,-1461.9,-2371.3,-2279.4,-16280.,-128.39,-19816.,-6318.9,-4265.5,-2677.4,76.164,2713.3,2474.1,2098.2,385.53,4665.4,1686.6,0.0000,7632.3,4449.7,4252.8,3658.0,0.0000,-431.10,-134.42,-110.97,-50.776,-143.60,-587.69,0.0000,-1071.6,-1568.8,-753.04,-1253.7
893.0000000000,104.13,2295.0,2365.1,1980.9,349.71,4214.7,970.97,23.913,6380.2,2689.4,3357.7,2001.5,0.0000,-7122.8,-7124.5,-1464.2,-2370.7,-2285.5,-16279.,-128.30,-19816.,-6318.5,-4264.8,-2676.6,75.762,2699.0,2461.0,2095.2,383.63,4662.2,1686.6,0.0000,7630.4,4449.7,4252.8,3658.0,0.0000,-428.89,-133.75,-110.66,-50.508,-143.68,-587.69,0.0000,-1071.6,-1568.7,-753.03,-1253.6
894.0000000000,103.73,2285.2,2357.2,1979.4,348.22,4224.6,970.95,22.432,6381.3,2690.5,3357.5,2001.8,0.0000,-7125.2,-7124.7,-1466.3,-2370.1,-2291.3,-16277.,-128.21,-19817.,-6318.2,-4264.2,-2675.7,75.458,2688.2,2451.2,2093.9,382.22,4662.1,1686.6,0.0000,7630.4,4449.7,4252.8,3658.0,0.0000,-427.24,-133.25,-110.46,-50.306,-143.86,-587.69,0.0000,-1071.6,-1568.6,-753.01,-1253.4
895.0000000000,103.43,2281.8,2353.0,1978.4,347.82,4233.1,970.95,22.558,6382.3,2690.0,3357.1,2002.1,0.0000,-7127.6,-7124.8,-1468.4,-2369.5,-2296.8,-16276.,-128.13,-19817.,-6317.8,-4263.6,-2674.8,213.95,2867.4,2614.9,2176.5,429.08,4754.0,1686.6,210.78,7710.1,4503.1,4302.4,3705.1,0.0000,-431.46,-137.51,-111.39,-51.032,-145.44,-587.69,-9.6410,-1072.6,-1568.5,-753.26,-1254.7
896.0000000000,103.64,2288.0,2356.2,1981.1,348.79,4244.9,970.95,19.737,6384.2,2688.1,3357.3,2002.1,0.0000,-7130.5,-7125.3,-1470.5,-2369.1,-2302.3,-16274.,-128.04,-19817.,-6317.5,-4262.9,-2674.0,76.310,2718.5,2478.8,2111.4,386.42,4698.0,1686.6,0.0000,7652.0,4449.8,4252.9,3658.1,0.0000,-432.19,-134.82,-111.49,-50.873,-145.34,-587.69,0.0000,-1071.8,-1568.4,-752.98,-1253.1
897.0000000000,103.69,2292.6,2361.7,1985.0,349.68,4262.4,970.95,19.736,6393.8,2687.0,3357.5,2002.3,0.0000,-7133.8,-7126.1,-1472.7,-2368.6,-2307.7,-16273.,-127.96,-19819.,-6317.1,-4262.3,-2673.1,224.69,2730.9,2687.4,2117.6,467.38,4719.1,1686.6,0.0000,7659.4,4449.7,4267.2,3676.5,0.0000,-434.22,-139.69,-111.89,-51.594,-145.95,-587.69,0.0000,-1071.9,-1568.3,-753.04,-1253.5
898.0000000000,104.02,2297.6,2365.8,1989.6,351.00,4267.7,970.96,19.734,6404.6,2687.1,3357.3,2002.6,0.0000,-7137.3,-7127.1,-1474.8,-2368.2,-2312.9,-16271.,-127.87,-19821.,-6316.7,-4261.7,-2672.3,76.717,2733.0,2492.1,2118.3,388.41,4711.3,1686.6,0.0000,7660.1,4449.7,4252.8,3658.0,0.0000,-434.62,-135.62,-111.94,-51.145,-146.12,-587.69,0.0000,-1071.9,-1568.1,-752.95,-1252.8
899.0000000000,103.93,2298.2,2367.8,1992.5,351.27,4274.0,970.96,18.694,6407.0,2687.2,3357.2,2003.0,0.0000,-7140.5,-7127.9,-1477.0,-2367.8,-2318.0,-16270.,-127.79,-19822.,-6316.3,-4261.0,-2671.4,76.498,2725.2,2484.9,2114.6,387.34,4704.2,1686.6,0.0000,7655.8,4449.7,4252.8,3658.0,0.0000,-433.44,-135.27,-111.70,-50.998,-146.07,-587.69,0.0000,-1071.9,-1568.0,-752.94,-1252.6
900.0000000000,103.91,2294.5,2364.3,1993.6,350.88,4287.5,970.96,16.087,6417.7,2687.3,3357.0,2003.0,0.0000,-7143.3,-7128.4,-1479.0,-2367.3,-2322.8,-16269.,-127.70,-19823.,-6315.9,-4260.4,-2670.6,76.199,2714.5,2475.2,2109.7,385.89,4695.0,1686.6,0.0000,7650.3,4449.7,4252.8,3658.0,0.0000,-431.80,-134.77,-111.38,-50.799,-145.95,-587.69,0.0000,-1071.9,-1567.9,-752.92,-1252.5
901.0000000000,103.77,2290.9,2362.9,1992.3,350.42,4289.7,970.96,14.256,6421.6,2688.0,3357.0,2003.0,0.0000,-7145.6,-7128.7,-1480.8,-2366.8,-2327.3,-16267.,-127.62,-19823.,-6315.4,-4259.8,-2669.7,159.67,2835.9,2577.7,2155.1,407.26,4717.0,1686.6,168.14,7682.3,4502.0,4278.4,3701.0,0.0000,-433.31,-137.23,-111.60,-51.073,-146.36,-587.69,-7.6905,-1072.4,-1567.8,-753.04,-1253.6
902.0000000000,103.57,2290.9,2364.9,1990.9,350.27,4291.9,970.96,12.440,6424.3,2688.3,3357.0,2003.0,0.0000,-7148.1,-7129.0,-1482.6,-2366.3,-2331.6,-16266.,-127.53,-19824.,-6315.0,-4259.2,-2668.8,76.303,2718.2,2478.6,2108.8,386.35,4691.4,1686.6,0.0000,7648.1,4449.7,4252.8,3658.0,0.0000,-432.50,-135.01,-111.40,-50.868,-146.17,-587.69,0.0000,-1071.9,-1567.7,-752.89,-1252.2
903.0000000000,103.35,2288.1,2363.5,1989.9,349.69,4291.6,970.96,12.440,6432.4,2688.4,3357.0,2003.1,0.0000,-7150.3,-7129.0,-1484.2,-2365.7,-2335.8,-16264.,-127.45,-19824.,-6314.6,-4258.5,-2668.0,76.023,2708.3,2469.5,2103.3,384.97,4680.3,1686.6,0.0000,7641.4,4449.7,4252.8,3658.0,0.0000,-430.95,-134.54,-111.07,-50.682,-145.97,-587.69,0.0000,-1071.9,-1567.6,-752.87,-1252.0
904.0000000000,103.20,2283.4,2359.0,1988.0,349.17,4288.6,970.97,12.439,6441.2,2688.5,3357.1,2003.1,0.0000,-7152.1,-7128.9,-1485.6,-2365.1,-2339.7,-16263.,-127.36,-19824.,-6314.2,-4257.9,-2667.1,131.28,2705.6,2467.1,2099.3,384.56,4670.8,1686.6,0.0000,7635.6,4449.7,4252.8,3658.0,0.0000,-430.57,-134.43,-110.90,-50.632,-145.83,-587.69,0.0000,-1071.9,-1567.5,-752.86,-1251.9
905.0000000000,102.86,2279.3,2356.3,1985.5,348.43,4283.3,970.97,11.673,6445.5,2689.1,3357.3,2003.1,0.0000,-7153.7,-7128.5,-1486.9,-2364.5,-2343.4,-16261.,-127.28,-19824.,-6313.8,-4257.3,-2666.3,75.651,2695.0,2457.4,2093.3,383.09,4658.4,1686.6,0.0000,7628.1,4449.7,4252.8,3658.0,0.0000,-428.92,-133.92,-110.54,-50.434,-145.58,-587.69,0.0000,-1071.8,-1567.3,-752.84,-1251.7
906.0000000000,102.59,2272.5,2350.7,1981.9,347.28,4276.6,970.97,8.7927,6444.3,2689.6,3357.3,2003.2,0.0000,-7154.7,-7128.0,-1488.1,-2363.9,-2346.8,-16260.,-127.19,-19824.,-6313.4,-4256.7,-2665.4,75.325,2683.4,2446.8,2086.8,381.48,4645.3,1686.6,0.0000,7620.2,4449.7,4252.8,3658.0,0.0000,-427.10,-133.35,-110.15,-50.217,-145.32,-587.69,0.0000,-1071.8,-1567.2,-752.83,-1251.6
907.0000000000,102.28,2264.5,2342.0,1977.4,346.08,4270.5,970.97,8.7931,6441.4,2689.1,3357.3,2003.4,0.0000,-7155.1,-7127.2,-1489.2,-2363.2,-2350.1,-16259.,-127.10,-19824.,-6313.0,-4256.1,-2664.5,74.983,2671.2,2435.7,2082.9,379.85,4639.0,1686.6,0.0000,7616.5,4449.7,4252.8,3658.0,0.0000,-425.18,-132.75,-109.84,-49.989,-145.26,-587.69,0.0000,-1071.8,-1567.1,-752.81,-1251.4
908.0000000000,101.77,2260.0,2337.9,1977.2,345.48,4264.9,970.97,8.7900,6437.9,2688.7,3357.3,2003.6,0.0000,-7155.4,-7126.4,-1490.2,-2362.5,-2353.3,-16257.,-127.02,-19824.,-6312.6,-4255.5,-2663.7,197.12,2772.0,2536.1,2114.2,410.43,4658.2,1686.6,100.96,7642.5,4491.4,4273.8,3692.0,0.0000,-428.16,-135.44,-110.18,-50.495,-145.52,-587.69,-4.6173,-1072.2,-1567.0,-752.91,-1252.3
909.0000000000,101.94,2269.8,2344.7,1978.1,346.91,4260.6,970.97,8.7965,6434.5,2688.3,3357.3,2003.7,0.0000,-7156.6,-7126.2,-1491.2,-2361.9,-2356.4,-16256.,-126.93,-19824.,-6312.2,-4254.9,-2662.8,373.50,2929.5,2773.0,2157.4,454.41,4702.5,1686.6,15.317,7656.0,4454.8,4307.2,3698.6,0.0000,-434.54,-141.68,-111.07,-51.456,-146.22,-587.69,-0.70051,-1072.3,-1566.9,-753.06,-1252.4
910.0000000000,102.53,2286.9,2359.1,1978.5,349.18,4258.5,970.97,8.8035,6431.4,2688.4,3357.5,2003.8,0.0000,-7159.1,-7126.8,-1492.3,-2361.4,-2359.5,-16254.,-126.85,-19823.,-6311.8,-4254.3,-2662.0,76.933,2740.7,2499.0,2092.7,388.96,4642.5,1686.6,0.0000,7618.2,4449.7,4252.8,3658.0,0.0000,-436.33,-136.26,-111.18,-51.288,-145.76,-587.69,0.0000,-1071.9,-1566.8,-752.76,-1251.0
911.0000000000,103.04,2297.0,2368.4,1979.2,350.74,4254.9,970.97,8.8037,6428.1,2688.5,3357.6,2003.6,0.0000,-7161.9,-7127.6,-1493.5,-2361.0,-2362.6,-16253.,-126.77,-19823.,-6311.4,-4253.7,-2661.1,76.824,2736.8,2495.5,2090.8,388.43,4638.8,1686.6,0.0000,7615.9,4449.7,4252.8,3658.0,0.0000,-435.76,-136.09,-111.06,-51.216,-145.78,-587.69,0.0000,-1071.9,-1566.6,-752.75,-1250.8
912.0000000000,103.36,2299.3,2370.9,1979.3,351.58,4250.7,970.94,8.8086,6425.1,2688.6,3357.6,2003.8,0.0000,-7164.5,-7128.2,-1494.5,-2360.5,-2365.4,-16251.,-126.68,-19822.,-6310.9,-4253.1,-2660.3,76.837,2737.3,2495.9,2090.1,388.48,4636.9,1686.6,0.0000,7614.8,4449.7,4252.8,3658.0,0.0000,-435.87,-136.14,-111.04,-51.225,-145.85,-587.69,0.0000,-1071.9,-1566.5,-752.73,-1250.7
913.0000000000,103.49,2298.9,2370.4,1985.4,351.52,4247.0,970.91,8.8092,6423.6,2689.1,3357.5,2003.9,0.0000,-7166.7,-7128.6,-1495.6,-2360.0,-2368.2,-16250.,-126.60,-19822.,-6310.5,-4252.5,-2659.4,76.568,2727.7,2487.2,2087.9,387.21,4633.9,1686.6,0.0000,7613.1,4449.7,4252.8,3658.0,0.0000,-434.39,-135.69,-110.82,-51.045,-145.88,-587.69,0.0000,-1071.9,-1566.4,-752.72,-1250.5
914.0000000000,103.31,2295.4,2366.6,1984.7,350.68,4244.4,970.89,8.8008,6423.3,2689.4,3357.4,2004.1,0.0000,-7168.3,-7128.8,-1496.6,-2359.5,-2370.9,-16249.,-126.51,-19821.,-6310.1,-4251.9,-2658.6,76.266,2716.9,2477.4,2085.4,385.77,4630.9,1686.6,0.0000,7611.3,4449.7,4252.8,3658.0,0.0000,-432.71,-135.17,-110.58,-50.844,-145.91,-587.69,0.0000,-1071.9,-1566.3,-752.70,-1250.4
915.0000000000,103.10,2289.1,2361.3,1983.0,349.67,4243.2,970.89,7.3176,6423.2,2690.2,3357.4,2004.2,0.0000,-7169.4,-7128.6,-1497.4,-2358.8,-2373.4,-16247.,-126.43,-19821.,-6309.7,-4251.3,-2657.7,75.937,2705.2,2466.7,2082.7,384.22,4627.8,1686.6,0.0000,7609.4,4449.7,4252.8,3658.0,0.0000,-430.87,-134.60,-110.32,-50.625,-145.94,-587.69,0.0000,-1071.9,-1566.2,-752.69,-1250.2
916.0000000000,102.80,2281.9,2354.9,1981.3,348.43,4244.4,970.89,7.3179,6421.7,2690.2,3357.5,2004.4,0.0000,-7170.0,-7128.1,-1498.3,-2358.1,-2375.9,-16246.,-126.34,-19820.,-6309.2,-4250.7,-2656.9,75.598,2693.1,2455.7,2080.0,382.62,4624.5,1686.6,0.0000,7607.5,4449.7,4252.8,3658.0,0.0000,-428.97,-134.01,-110.06,-50.399,-145.96,-587.69,0.0000,-1071.9,-1566.1,-752.67,-1250.1
917.0000000000,102.62,2273.5,2347.0,1979.9,347.07,4244.7,970.89,7.3182,6419.8,2690.0,3357.7,2004.6,0.0000,-7170.0,-7127.3,-1499.0,-2357.4,-2378.3,-16244.,-126.26,-19819.,-6308.8,-4250.1,-2656.0,75.251,2680.8,2444.4,2077.2,380.98,4621.2,1686.6,0.0000,7605.6,4449.7,4252.8,3658.0,0.0000,-427.01,-133.39,-109.78,-50.168,-145.98,-587.69,0.0000,-1071.9,-1566.0,-752.66,-1249.9
918.0000000000,102.30,2264.8,2338.0,1978.2,345.62,4241.4,970.90,7.3239,6418.0,2690.3,3357.7,2004.6,0.0000,-7169.4,-7126.3,-1499.8,-2356.6,-2380.6,-16243.,-126.18,-19819.,-6308.4,-4249.5,-2655.2,74.895,2668.1,2432.8,2074.4,379.29,4617.8,1686.6,0.0000,7603.6,4449.7,4252.8,3658.0,0.0000,-424.99,-132.76,-109.50,-49.930,-145.99,-587.69,0.0000,-1071.9,-1565.8,-752.64,-1249.8
919.0000000000,101.98,2261.8,2333.7,1976.3,345.05,4238.7,970.90,7.3353,6416.2,2690.1,3357.7,2004.6,0.0000,-7168.8,-7125.3,-1500.5,-2355.9,-2382.8,-16241.,-126.09,-19818.,-6307.9,-4248.9,-2654.3,228.69,2749.0,2501.5,2096.8,400.02,4639.4,1686.6,4.4722,7615.3,4453.0,4266.5,3667.4,0.0000,-428.42,-134.85,-109.89,-50.431,-146.22,-587.69,-0.20452,-1072.1,-1565.7,-752.70,-1249.9
920.0000000000,102.14,2265.0,2336.2,1975.0,345.50,4236.4,970.90,7.3356,6414.5,2689.1,3357.6,2004.7,0.0000,-7168.6,-7124.7,-1501.2,-2355.2,-2384.9,-16240.,-126.01,-19817.,-6307.5,-4248.4,-2653.5,75.416,2686.6,2449.8,2075.6,381.71,4615.1,1686.6,0.0000,7601.9,4449.7,4252.8,3658.0,0.0000,-427.96,-133.68,-109.81,-50.277,-146.12,-587.69,0.0000,-1071.9,-1565.6,-752.61,-1249.5
921.0000000000,102.03,2264.5,2336.4,1974.4,345.25,4234.2,970.90,7.0935,6412.8,2689.0,3357.5,2004.8,0.0000,-7168.4,-7124.1,-1501.9,-2354.5,-2386.9,-16238.,-125.93,-19817.,-6307.0,-4247.8,-2652.6,75.221,2679.7,2443.4,2073.4,380.77,4611.7,1686.6,0.0000,7599.8,4449.7,4252.8,3658.0,0.0000,-426.86,-133.33,-109.64,-50.147,-146.13,-587.69,0.0000,-1071.9,-1565.5,-752.60,-1249.3
922.0000000000,102.05,2260.8,2333.0,1973.3,345.08,4231.2,970.90,5.8434,6412.1,2689.0,3357.4,2004.8,0.0000,-7168.0,-7123.4,-1502.5,-2353.8,-2388.9,-16237.,-125.85,-19816.,-6306.5,-4247.2,-2651.8,74.965,2670.6,2435.1,2071.0,379.56,4608.3,1686.6,0.0000,7597.8,4449.7,4252.8,3658.0,0.0000,-425.40,-132.87,-109.42,-49.976,-146.13,-587.69,0.0000,-1071.9,-1565.4,-752.58,-1249.2
923.0000000000,101.89,2254.5,2327.7,1971.4,344.18,4228.2,970.90,5.8438,6416.9,2689.3,3357.5,2004.9,0.0000,-7167.2,-7122.4,-1503.2,-2353.0,-2390.8,-16235.,-125.76,-19815.,-6306.0,-4246.6,-2650.9,74.675,2660.2,2425.7,2068.4,378.18,4604.7,1686.6,0.0000,7595.7,4449.7,4252.8,3658.0,0.0000,-423.75,-132.35,-109.18,-49.783,-146.12,-587.69,0.0000,-1071.9,-1565.3,-752.57,-1249.0
924.0000000000,101.63,2247.4,2319.8,1970.1,343.08,4225.2,970.90,5.8441,6415.2,2689.2,3357.6,2005.0,0.0000,-7166.0,-7121.3,-1503.7,-2352.2,-2392.6,-16234.,-125.68,-19814.,-6305.5,-4246.0,-2650.1,74.361,2649.1,2415.5,2066.5,376.71,4603.3,1686.6,0.0000,7594.9,4449.7,4252.8,3658.0,0.0000,-421.96,-131.78,-108.96,-49.574,-146.18,-587.69,0.0000,-1071.9,-1565.2,-752.55,-1248.9
925.0000000000,101.53,2239.1,2311.9,1975.4,341.95,4222.7,970.90,6.6895,6413.7,2688.9,3357.5,2005.2,0.0000,-7164.3,-7119.9,-1504.2,-2351.4,-2394.3,-16232.,-125.60,-19813.,-6305.1,-4245.4,-2649.3,74.036,2637.5,2405.0,2064.8,375.19,4602.7,1686.6,0.0000,7594.6,4449.7,4252.8,3658.0,0.0000,-420.10,-131.19,-108.73,-49.358,-146.27,-587.69,0.0000,-1071.9,-1565.0,-752.54,-1248.8
926.0000000000,101.25,2230.5,2303.8,1973.9,340.67,4220.6,970.90,6.6197,6412.5,2688.7,3357.4,2005.4,0.0000,-7162.3,-7118.4,-1504.7,-2350.5,-2396.0,-16231.,-125.52,-19812.,-6304.6,-4244.8,-2648.4,73.706,2625.7,2394.2,2063.2,373.65,4602.1,1686.6,0.0000,7594.3,4449.7,4252.8,3658.0,0.0000,-418.20,-130.58,-108.51,-49.137,-146.35,-587.69,0.0000,-1071.9,-1564.9,-752.52,-1248.6
927.0000000000,101.11,2222.0,2294.9,1972.8,339.36,4218.4,970.91,6.2661,6411.4,2688.7,3357.3,2005.6,0.0000,-7159.9,-7116.7,-1505.2,-2349.6,-2397.7,-16229.,-125.44,-19811.,-6304.1,-4244.3,-2647.6,73.372,2613.9,2383.4,2061.5,372.09,4601.6,1686.6,0.0000,7594.0,4449.7,4252.8,3658.0,0.0000,-416.28,-129.96,-108.28,-48.915,-146.44,-587.69,0.0000,-1071.9,-1564.8,-752.51,-1248.5
928.0000000000,100.77,2212.9,2285.3,1972.0,338.08,4216.3,970.91,6.2665,6410.2,2688.7,3357.6,2005.8,0.0000,-7157.1,-7114.8,-1505.6,-2348.7,-2399.3,-16228.,-125.37,-19810.,-6303.6,-4243.7,-2646.7,73.036,2601.9,2372.5,2059.8,370.52,4601.0,1686.6,0.0000,7593.7,4449.7,4252.8,3658.0,0.0000,-414.34,-129.33,-108.05,-48.691,-146.52,-587.69,0.0000,-1071.9,-1564.7,-752.49,-1248.3
929.0000000000,100.38,2204.1,2275.9,1970.9,336.73,4214.6,970.91,6.2669,6409.1,2688.9,3357.7,2005.9,0.0000,-7153.8,-7112.7,-1506.1,-2347.7,-2400.9,-16226.,-125.29,-19810.,-6303.1,-4243.1,-2645.9,72.698,2589.8,2361.5,2058.1,368.93,4600.4,1686.6,0.0000,7593.4,4449.7,4252.8,3658.0,0.0000,-412.38,-128.70,-107.82,-48.465,-146.60,-587.69,0.0000,-1072.0,-1564.6,-752.48,-1248.2
930.0000000000,99.921,2194.6,2267.2,1969.5,335.35,4213.4,970.90,6.2672,6408.2,2689.0,3357.5,2006.0,0.0000,-7150.3,-7110.5,-1506.5,-2346.7,-2402.5,-16225.,-125.21,-19809.,-6302.7,-4242.5,-2645.1,72.355,2577.6,2350.4,2056.4,367.33,4599.8,1686.6,0.0000,7593.1,4449.7,4252.8,3658.0,0.0000,-410.39,-128.05,-107.58,-48.237,-146.68,-587.69,0.0000,-1072.0,-1564.5,-752.47,-1248.0
931.0000000000,99.576,2185.1,2258.0,1968.1,333.93,4219.7,970.89,6.2676,6407.4,2689.3,3357.4,2006.0,0.0000,-7146.5,-7108.2,-1506.9,-2345.7,-2404.0,-16223.,-125.14,-19808.,-6302.2,-4241.9,-2644.2,72.018,2565.6,2339.4,2054.7,365.75,4599.2,1686.6,0.0000,7592.8,4449.7,4252.8,3658.0,0.0000,-408.42,-127.41,-107.35,-48.012,-146.75,-587.69,0.0000,-1072.0,-1564.4,-752.45,-1247.9
932.0000000000,99.233,2175.4,2248.6,1966.7,332.57,4218.6,970.89,6.2680,6406.8,2689.6,3357.4,2006.2,0.0000,-7142.3,-7105.8,-1507.3,-2344.7,-2405.5,-16222.,-125.06,-19807.,-6301.7,-4241.4,-2643.4,71.680,2553.6,2328.4,2053.0,364.17,4598.6,1686.6,0.0000,7592.5,4449.7,4252.8,3658.0,0.0000,-406.45,-126.77,-107.12,-47.787,-146.83,-587.69,0.0000,-1072.0,-1564.3,-752.44,-1247.7
933.0000000000,98.890,2165.7,2239.4,1965.5,331.20,4217.5,970.89,5.0553,6406.2,2690.2,3357.4,2006.5,0.0000,-7138.0,-7103.3,-1507.6,-2343.6,-2407.0,-16220.,-124.99,-19806.,-6301.2,-4240.8,-2642.5,71.345,2541.6,2317.5,2051.4,362.61,4598.1,1686.6,0.0000,7592.3,4449.7,4252.8,3658.0,0.0000,-404.49,-126.13,-106.89,-47.563,-146.91,-587.69,0.0000,-1072.0,-1564.1,-752.42,-1247.6
934.0000000000,98.549,2156.2,2230.5,1964.3,329.90,4216.5,970.89,5.0372,6405.6,2690.3,3357.5,2006.5,0.0000,-7133.4,-7100.6,-1507.9,-2342.5,-2408.4,-16219.,-124.92,-19805.,-6300.8,-4240.2,-2641.7,71.012,2529.8,2306.7,2049.9,361.05,4597.9,1686.6,0.0000,7592.3,4449.7,4252.8,3658.0,0.0000,-402.54,-125.49,-106.67,-47.341,-146.99,-587.69,0.0000,-1072.0,-1564.0,-752.41,-1247.4
935.0000000000,98.197,2146.7,2220.8,1962.9,328.55,4220.9,970.86,5.1704,6405.1,2690.5,3357.6,2006.6,0.0000,-7128.5,-7097.9,-1508.3,-2341.5,-2409.7,-16217.,-124.84,-19804.,-6300.3,-4239.6,-2640.9,70.684,2518.1,2296.1,2048.4,359.52,4597.8,1686.6,0.0000,7592.3,4449.7,4252.8,3658.0,0.0000,-400.61,-124.86,-106.45,-47.123,-147.08,-587.69,0.0000,-1072.0,-1563.9,-752.39,-1247.3
936.0000000000,97.718,2137.1,2211.1,1961.8,327.17,4222.8,970.85,5.1708,6404.6,2690.6,3357.5,2006.8,0.0000,-7123.4,-7095.1,-1508.6,-2340.3,-2411.1,-16216.,-124.77,-19802.,-6299.8,-4239.0,-2640.0,70.362,2506.6,2285.6,2046.9,358.02,4597.7,1686.6,0.0000,7592.3,4449.7,4252.8,3658.0,0.0000,-398.70,-124.23,-106.23,-46.908,-147.16,-587.69,0.0000,-1072.0,-1563.8,-752.38,-1247.2
937.0000000000,97.387,2127.7,2201.2,1960.5,325.79,4222.2,970.83,5.1713,6404.1,2690.3,3357.4,2006.9,0.0000,-7118.0,-7092.1,-1508.8,-2339.2,-2412.4,-16214.,-124.69,-19801.,-6299.4,-4238.5,-2639.2,70.036,2495.0,2275.0,2045.5,356.50,4597.5,1686.6,0.0000,7592.2,4449.7,4252.8,3658.0,0.0000,-396.78,-123.60,-106.02,-46.690,-147.24,-587.69,0.0000,-1072.0,-1563.7,-752.37,-1247.0
938.0000000000,97.056,2118.3,2191.3,1959.1,324.49,4221.7,970.80,4.1896,6403.7,2690.4,3357.4,2007.0,0.0000,-7112.5,-7089.1,-1509.1,-2338.1,-2413.7,-16213.,-124.62,-19800.,-6298.9,-4237.9,-2638.4,69.709,2483.4,2264.4,2044.0,354.97,4597.4,1686.6,0.0000,7592.2,4449.7,4252.8,3658.0,0.0000,-394.85,-122.96,-105.80,-46.473,-147.32,-587.69,0.0000,-1072.1,-1563.6,-752.35,-1246.9
939.0000000000,96.726,2108.8,2181.8,1957.9,323.19,4221.0,970.81,3.6780,6403.3,2690.5,3357.5,2007.1,0.0000,-7106.7,-7086.2,-1509.4,-2336.9,-2414.9,-16211.,-124.54,-19799.,-6298.5,-4237.3,-2637.5,69.390,2472.0,2254.0,2042.5,353.48,4597.2,1686.6,0.0000,7592.2,4449.7,4252.8,3658.0,0.0000,-392.95,-122.33,-105.58,-46.260,-147.40,-587.69,0.0000,-1072.1,-1563.5,-752.34,-1246.7
940.0000000000,96.399,2099.1,2172.4,1956.6,321.91,4220.5,970.80,3.6785,6403.2,2690.6,3357.6,2007.2,0.0000,-7100.7,-7083.1,-1509.6,-2335.8,-2416.1,-16210.,-124.47,-19798.,-6298.0,-4236.7,-2636.7,69.078,2460.9,2243.9,2041.1,352.03,4597.1,1686.6,0.0000,7592.2,4449.7,4252.8,3658.0,0.0000,-391.10,-121.72,-105.38,-46.052,-147.47,-587.69,0.0000,-1072.1,-1563.4,-752.32,-1246.6
941.0000000000,95.860,2090.2,2163.2,1955.3,320.64,4220.0,970.76,3.7799,6403.1,2690.7,3357.5,2007.4,0.0000,-7094.5,-7080.0,-1509.8,-2334.6,-2417.3,-16208.,-124.40,-19797.,-6297.6,-4236.2,-2635.8,68.769,2449.9,2233.9,2039.7,350.59,4597.0,1686.6,0.0000,7592.2,4449.7,4252.8,3658.0,0.0000,-389.26,-121.11,-105.17,-45.846,-147.55,-587.69,0.0000,-1072.1,-1563.3,-752.31,-1246.4
942.0000000000,95.369,2081.3,2154.0,1954.1,319.39,4219.6,970.76,3.7838,6402.9,2690.8,3357.6,2007.5,0.0000,-7088.2,-7076.8,-1510.0,-2333.4,-2418.5,-16207.,-124.32,-19796.,-6297.1,-4235.6,-2635.0,68.468,2439.1,2224.1,2038.4,349.18,4596.8,1686.6,0.0000,7592.2,4449.7,4252.8,3658.0,0.0000,-387.46,-120.51,-104.97,-45.645,-147.62,-587.69,0.0000,-1072.1,-1563.2,-752.29,-1246.3
943.0000000000,95.009,2073.9,2146.1,1953.0,318.43,4219.1,970.77,3.7843,6402.7,2690.9,3357.7,2007.7,0.0000,-7081.9,-7073.6,-1510.2,-2332.2,-2419.7,-16205.,-124.25,-19795.,-6296.7,-4235.0,-2634.2,69.089,2442.5,2224.1,2038.4,349.18,4596.8,1686.6,0.0000,7592.2,4449.7,4252.8,3658.0,0.0000,-387.37,-120.44,-104.97,-45.646,-147.69,-587.69,0.0000,-1072.1,-1563.0,-752.28,-1246.1
944.0000000000,94.863,2069.6,2140.9,1952.0,317.93,4218.7,970.77,3.7848,6402.6,2691.0,3357.6,2007.8,0.0000,-7075.8,-7070.6,-1510.4,-2331.0,-2420.8,-16204.,-124.18,-19794.,-6296.2,-4234.4,-2633.3,68.369,2435.6,2220.9,2037.9,348.72,4596.8,1686.6,0.0000,7592.2,4449.7,4252.8,3658.0,0.0000,-386.71,-120.20,-104.90,-45.579,-147.76,-587.69,0.0000,-1072.1,-1562.9,-752.27,-1246.0
945.0000000000,94.701,2064.8,2136.0,1951.2,317.26,4218.4,970.77,3.7853,6402.4,2691.1,3357.7,2007.9,0.0000,-7069.7,-7067.6,-1510.6,-2329.9,-2421.9,-16202.,-124.10,-19793.,-6295.7,-4233.9,-2632.5,68.093,2425.8,2211.9,2036.7,347.43,4596.7,1686.6,0.0000,7592.2,4449.7,4252.8,3658.0,0.0000,-385.06,-119.65,-104.72,-45.396,-147.83,-587.69,0.0000,-1072.1,-1562.8,-752.25,-1245.9
946.0000000000,94.497,2058.0,2129.2,1950.4,316.45,4218.0,970.77,3.7858,6402.3,2691.0,3357.7,2008.1,0.0000,-7063.6,-7064.6,-1510.8,-2328.7,-2422.9,-16201.,-124.03,-19792.,-6295.3,-4233.3,-2631.7,67.810,2415.7,2202.7,2035.4,346.11,4596.6,1686.6,0.0000,7592.1,4449.7,4252.8,3658.0,0.0000,-383.36,-119.09,-104.53,-45.207,-147.90,-587.69,0.0000,-1072.1,-1562.7,-752.24,-1245.7
947.0000000000,94.283,2050.2,2121.2,1949.5,315.46,4217.8,970.77,3.7428,6402.2,2691.1,3357.7,2008.2,0.0000,-7057.3,-7061.5,-1510.9,-2327.5,-2424.0,-16199.,-123.96,-19791.,-6294.8,-4232.7,-2630.8,67.522,2405.4,2193.3,2034.1,344.76,4596.5,1686.6,0.0000,7592.1,4449.7,4252.8,3658.0,0.0000,-381.63,-118.51,-104.34,-45.014,-147.96,-587.69,0.0000,-1072.1,-1562.6,-752.22,-1245.6
948.0000000000,94.016,2042.1,2112.8,1948.4,314.27,4217.5,970.77,3.6753,6402.1,2691.2,3357.6,2008.4,0.0000,-7050.9,-7058.4,-1511.1,-2326.3,-2425.0,-16198.,-123.88,-19790.,-6294.4,-4232.1,-2630.0,67.231,2395.1,2183.9,2032.9,343.41,4596.4,1686.6,0.0000,7592.1,4449.7,4252.8,3658.0,0.0000,-379.89,-117.93,-104.14,-44.821,-148.02,-587.69,0.0000,-1072.2,-1562.5,-752.21,-1245.4
949.0000000000,93.725,2033.8,2104.3,1947.3,313.10,4217.2,970.77,3.7272,6401.9,2691.1,3357.6,2008.5,0.0000,-7044.3,-7055.2,-1511.2,-2325.1,-2426.0,-16196.,-123.81,-19789.,-6293.9,-4231.6,-2629.2,66.944,2384.8,2174.6,2031.6,342.07,4596.3,1686.6,0.0000,7592.1,4449.7,4252.8,3658.0,0.0000,-378.16,-117.36,-103.95,-44.629,-148.09,-587.69,0.0000,-1072.2,-1562.4,-752.20,-1245.3
950.0000000000,93.433,2025.7,2095.9,1945.6,311.95,4215.7,970.77,3.2830,6401.5,2691.2,3357.6,2008.6,0.0000,-7037.5,-7052.0,-1511.3,-2323.9,-2426.9,-16195.,-123.74,-19788.,-6293.5,-4231.0,-2628.3,66.659,2374.7,2165.3,2019.3,340.55,4567.7,1686.6,0.0000,7574.8,4449.7,4252.8,3658.0,0.0000,-376.45,-116.79,-103.39,-44.439,-147.20,-587.69,0.0000,-1072.0,-1562.3,-752.18,-1245.1
951.0000000000,93.142,2017.8,2087.3,1941.0,310.71,4208.5,970.74,2.2369,6399.8,2691.3,3357.6,2008.8,0.0000,-7030.6,-7048.7,-1511.1,-2322.6,-2427.6,-16193.,-123.66,-19786.,-6293.0,-4230.4,-2627.5,66.377,2364.7,2156.2,2004.5,339.00,4532.4,1686.6,0.0000,7553.4,4449.7,4252.8,3658.0,0.0000,-374.76,-116.22,-102.73,-44.251,-146.10,-587.69,0.0000,-1071.9,-1562.2,-752.17,-1245.0
952.0000000000,92.853,2009.7,2078.8,1933.3,309.43,4195.7,970.72,2.2512,6396.1,2691.2,3357.6,2008.9,0.0000,-7023.6,-7045.4,-1510.8,-2321.4,-2428.0,-16191.,-123.59,-19785.,-6292.5,-4229.8,-2626.7,66.099,2354.7,2147.1,1989.9,337.47,4497.6,1686.6,0.0000,7532.3,4449.7,4252.8,3658.0,0.0000,-373.08,-115.66,-102.09,-44.066,-145.00,-587.69,0.0000,-1071.7,-1562.1,-752.15,-1244.8
953.0000000000,92.567,2001.7,2070.3,1923.0,308.09,4179.7,970.69,2.5954,6391.1,2691.2,3357.6,2009.0,0.0000,-7016.5,-7042.1,-1510.2,-2320.1,-2427.9,-16190.,-123.52,-19784.,-6292.1,-4229.3,-2625.9,65.826,2345.0,2138.3,1975.5,335.97,4463.2,1686.6,0.0000,7511.4,4449.7,4252.8,3658.0,0.0000,-371.43,-115.11,-101.46,-43.884,-143.90,-587.69,0.0000,-1071.6,-1562.0,-752.14,-1244.7
954.0000000000,92.267,1993.9,2061.7,1911.2,306.73,4161.6,970.67,2.6504,6384.5,2691.3,3357.6,2009.1,0.0000,-7009.3,-7038.7,-1509.4,-2318.9,-2427.5,-16188.,-123.45,-19783.,-6291.6,-4228.7,-2625.0,65.554,2335.3,2129.4,1961.1,334.48,4428.9,1686.6,0.0000,7490.6,4449.7,4252.8,3658.0,0.0000,-369.79,-114.56,-100.82,-43.702,-142.80,-587.69,0.0000,-1071.4,-1561.8,-752.12,-1244.6
955.0000000000,91.989,1986.7,2053.7,1898.9,305.49,4142.6,970.65,2.5643,6375.7,2691.2,3357.7,2009.2,0.0000,-7002.0,-7035.4,-1508.3,-2317.6,-2426.9,-16187.,-123.37,-19782.,-6291.1,-4228.1,-2624.2,65.444,2331.4,2125.9,1950.6,333.80,4402.9,1686.6,0.43388E-01,7474.8,4449.7,4252.8,3658.0,0.0000,-369.06,-114.30,-100.41,-43.630,-141.97,-587.69,-0.19837E-02,-1071.3,-1561.7,-752.11,-1244.4
956.0000000000,91.950,1980.9,2047.6,1887.3,304.56,4126.4,970.65,2.4871,6363.5,2691.4,3357.7,2009.3,0.0000,-6994.8,-7032.2,-1507.2,-2316.4,-2426.1,-16185.,-123.30,-19780.,-6290.7,-4227.6,-2623.4,65.237,2324.1,2119.1,1938.8,332.65,4374.6,1686.6,0.0000,7457.7,4449.7,4252.8,3658.0,0.0000,-367.78,-113.86,-99.899,-43.492,-141.05,-587.69,0.0000,-1071.2,-1561.6,-752.10,-1244.3
957.0000000000,91.594,1975.7,2042.2,1876.4,303.68,4106.6,970.65,2.4877,6349.4,2691.5,3357.7,2009.5,0.0000,-6987.7,-7029.0,-1505.9,-2315.1,-2425.3,-16183.,-123.23,-19779.,-6290.2,-4227.0,-2622.5,65.406,2323.7,2119.3,1931.1,332.83,4354.7,1686.6,0.0000,7445.6,4449.7,4252.9,3658.0,0.0000,-367.62,-113.79,-99.631,-43.487,-140.41,-587.69,0.0000,-1071.1,-1561.5,-752.08,-1244.1
958.0000000000,91.379,1976.3,2041.9,1866.4,303.85,4084.6,970.65,2.4290,6335.0,2691.6,3357.7,2009.6,0.0000,-6981.1,-7026.2,-1504.6,-2313.9,-2424.3,-16182.,-123.16,-19778.,-6289.7,-4226.4,-2621.7,70.393,2355.8,2148.5,1929.9,336.50,4342.0,1686.6,0.0000,7437.5,4449.7,4253.0,3658.0,0.0000,-371.82,-115.15,-99.963,-43.997,-139.98,-587.69,0.0000,-1071.0,-1561.4,-752.07,-1244.0
959.0000000000,91.623,1984.1,2047.6,1857.8,305.01,4064.3,970.65,2.2981,6321.1,2691.7,3357.7,2009.7,0.0000,-6975.5,-7023.9,-1503.4,-2312.9,-2423.3,-16180.,-123.09,-19776.,-6289.3,-4225.9,-2620.9,66.112,2355.2,2147.6,1917.9,336.30,4310.3,1686.6,0.0000,7418.4,4449.7,4252.8,3658.0,0.0000,-372.41,-115.20,-99.632,-44.075,-138.94,-587.69,0.0000,-1070.8,-1561.3,-752.05,-1243.8
960.0000000000,91.641,1988.2,2051.4,1849.8,305.33,4042.9,970.65,2.3139,6307.5,2691.7,3357.7,2009.8,0.0000,-6970.4,-7021.9,-1502.1,-2311.8,-2422.3,-16179.,-123.02,-19775.,-6288.8,-4225.3,-2620.1,66.037,2352.5,2145.1,1905.5,335.74,4279.0,1686.6,0.0000,7399.4,4449.7,4252.8,3658.0,0.0000,-371.90,-115.01,-99.168,-44.025,-137.91,-587.69,0.0000,-1070.7,-1561.2,-752.04,-1243.7
961.0000000000,91.580,1987.9,2051.0,1840.9,305.63,4019.9,970.66,2.5263,6294.0,2691.8,3357.7,2009.9,0.0000,-6965.3,-7019.9,-1500.8,-2310.8,-2420.9,-16177.,-122.94,-19773.,-6288.3,-4224.7,-2619.2,65.889,2347.3,2140.3,1892.7,334.85,4247.5,1686.6,0.0000,7380.3,4449.7,4252.8,3658.0,0.0000,-370.98,-114.70,-98.656,-43.926,-136.86,-587.69,0.0000,-1070.5,-1561.1,-752.03,-1243.6
962.0000000000,91.635,1987.2,2050.6,1830.9,305.56,3997.5,970.66,2.8007,6280.9,2691.9,3357.8,2010.0,0.0000,-6960.4,-7017.9,-1499.4,-2309.7,-2419.5,-16175.,-122.87,-19772.,-6287.9,-4224.1,-2618.4,66.178,2377.4,2173.9,1899.2,339.19,4253.2,1686.6,1.8844,7382.7,4450.3,4254.4,3658.5,0.0000,-372.56,-115.67,-98.886,-44.137,-136.96,-587.69,-0.86149E-01,-1070.5,-1561.0,-752.02,-1243.4
963.0000000000,91.768,1990.4,2052.9,1823.0,306.00,3979.5,970.66,2.8013,6269.7,2692.0,3357.8,2010.2,0.0000,-6955.8,-7016.1,-1498.0,-2308.7,-2418.0,-16174.,-122.80,-19770.,-6287.4,-4223.6,-2617.6,66.340,2375.8,2155.0,1897.1,336.86,4234.3,1686.6,3.6624,7375.1,4449.7,4252.8,3658.0,0.0000,-373.37,-115.38,-98.768,-44.226,-136.38,-587.69,-0.16743,-1070.5,-1560.9,-752.00,-1243.3
964.0000000000,91.848,1992.9,2055.4,1816.5,306.11,3963.9,970.66,2.8040,6259.4,2692.1,3357.8,2010.2,0.0000,-6951.5,-7014.5,-1496.6,-2307.7,-2416.5,-16172.,-122.73,-19769.,-6286.9,-4223.0,-2616.8,66.221,2359.1,2151.1,1877.8,336.11,4205.1,1686.6,0.0000,7354.4,4449.7,4252.8,3658.0,0.0000,-372.61,-115.13,-98.316,-44.147,-135.42,-587.69,0.0000,-1070.3,-1560.8,-751.98,-1243.1
965.0000000000,91.831,1991.6,2055.0,1809.5,305.90,3945.3,970.66,2.8075,6247.5,2692.2,3357.8,2010.4,0.0000,-6947.2,-7012.9,-1495.2,-2306.7,-2414.9,-16171.,-122.66,-19767.,-6286.5,-4222.4,-2615.9,66.032,2352.4,2145.0,1865.4,335.04,4175.0,1686.6,0.0000,7336.1,4449.7,4252.8,3658.0,0.0000,-371.47,-114.76,-97.795,-44.022,-134.41,-587.69,0.0000,-1070.2,-1560.7,-751.97,-1243.0
966.0000000000,91.781,1988.6,2052.6,1800.9,305.32,3923.4,970.66,2.8615,6234.3,2692.3,3357.8,2010.5,0.0000,-6942.8,-7011.1,-1493.7,-2305.7,-2413.1,-16169.,-122.59,-19766.,-6286.0,-4221.9,-2615.1,65.821,2344.8,2138.1,1853.0,333.85,4144.9,1686.6,0.0000,7317.9,4449.7,4252.8,3658.0,0.0000,-370.21,-114.34,-97.259,-43.881,-133.40,-587.69,0.0000,-1070.0,-1560.5,-751.95,-1242.9
967.0000000000,91.366,1983.9,2048.7,1791.5,304.39,3899.7,970.66,2.9147,6221.1,2692.5,3357.8,2010.6,0.0000,-6938.2,-7009.2,-1492.1,-2304.6,-2411.1,-16167.,-122.52,-19764.,-6285.5,-4221.3,-2614.3,65.596,2336.8,2130.8,1840.4,332.61,4114.9,1686.6,0.0000,7299.7,4449.7,4252.8,3658.0,0.0000,-368.87,-113.90,-96.714,-43.731,-132.39,-587.69,0.0000,-1069.8,-1560.4,-751.94,-1242.7
968.0000000000,91.090,1978.9,2043.6,1781.1,303.39,3877.6,970.66,2.7350,6209.6,2692.6,3357.8,2010.7,0.0000,-6933.3,-7007.3,-1490.4,-2303.6,-2408.8,-16166.,-122.45,-19762.,-6285.1,-4220.7,-2613.5,65.434,2331.1,2125.5,1830.8,331.70,4091.8,1686.6,0.0000,7285.7,4449.7,4252.8,3658.0,0.0000,-367.88,-113.57,-96.302,-43.623,-131.60,-587.69,0.0000,-1069.7,-1560.3,-751.93,-1242.6
969.0000000000,90.682,1975.5,2039.5,1770.6,302.60,3858.0,970.66,2.5614,6197.9,2692.7,3357.8,2010.9,0.0000,-6928.4,-7005.3,-1488.5,-2302.5,-2406.5,-16164.,-122.38,-19760.,-6284.6,-4220.2,-2612.7,67.066,2330.4,2124.9,1821.6,331.45,4068.1,1686.6,0.0000,7271.3,4449.7,4252.8,3658.0,0.0000,-367.70,-113.49,-95.977,-43.610,-130.78,-587.69,0.0000,-1069.6,-1560.2,-751.91,-1242.4
970.0000000000,90.515,1972.8,2036.8,1760.7,301.83,3837.3,970.65,2.5619,6184.9,2692.8,3357.8,2011.0,0.0000,-6923.5,-7003.3,-1486.7,-2301.4,-2404.0,-16162.,-122.31,-19759.,-6284.2,-4219.6,-2611.8,65.196,2322.6,2117.8,1809.6,330.24,4039.4,1686.6,0.0000,7253.8,4449.7,4252.8,3658.0,0.0000,-366.40,-113.06,-95.453,-43.464,-129.80,-587.69,0.0000,-1069.4,-1560.1,-751.90,-1242.3
971.0000000000,90.328,1968.4,2032.5,1751.2,300.91,3818.3,970.65,2.5625,6170.4,2693.0,3357.8,2011.1,0.0000,-6918.4,-7001.3,-1484.8,-2300.3,-2401.4,-16160.,-122.23,-19757.,-6283.7,-4219.0,-2611.0,64.975,2314.7,2110.6,1797.7,329.03,4011.0,1686.6,0.0000,7236.6,4449.7,4252.8,3658.0,0.0000,-365.09,-112.63,-94.932,-43.317,-128.82,-587.69,0.0000,-1069.3,-1560.0,-751.88,-1242.2
972.0000000000,90.147,1963.1,2026.8,1741.2,299.96,3797.4,970.66,2.5631,6155.2,2693.1,3357.8,2011.3,0.0000,-6913.2,-6999.2,-1482.8,-2299.2,-2398.7,-16159.,-122.16,-19755.,-6283.2,-4218.4,-2610.2,64.760,2307.0,2103.6,1786.1,327.84,3983.1,1686.6,0.0000,7219.7,4449.7,4252.8,3658.0,0.0000,-363.81,-112.21,-94.422,-43.173,-127.86,-587.69,0.0000,-1069.1,-1559.9,-751.87,-1242.0
973.0000000000,89.935,1957.8,2021.4,1730.7,298.93,3772.8,970.66,2.5636,6140.1,2693.2,3357.8,2011.5,0.0000,-6907.9,-6997.1,-1480.7,-2298.1,-2395.8,-16157.,-122.09,-19753.,-6282.8,-4217.9,-2609.4,64.612,2301.8,2098.8,1775.5,326.98,3957.4,1686.6,0.0000,7204.1,4449.7,4252.8,3658.0,0.0000,-362.90,-111.90,-93.986,-43.075,-126.97,-587.69,0.0000,-1069.0,-1559.8,-751.85,-1241.9
974.0000000000,89.656,1952.9,2016.0,1720.1,297.92,3749.0,970.66,2.4221,6126.0,2693.3,3357.8,2011.6,0.0000,-6902.4,-6994.9,-1478.6,-2297.0,-2392.8,-16155.,-122.02,-19751.,-6282.3,-4217.3,-2608.6,64.365,2293.0,2090.8,1763.3,325.64,3928.5,1686.6,0.0000,7186.6,4449.7,4252.8,3658.0,0.0000,-361.44,-111.42,-93.442,-42.910,-125.97,-587.69,0.0000,-1068.9,-1559.7,-751.84,-1241.7
975.0000000000,89.428,1946.9,2009.9,1709.7,296.83,3725.6,970.66,2.4001,6111.9,2693.4,3357.8,2011.8,0.0000,-6896.7,-6992.7,-1476.5,-2295.9,-2389.7,-16154.,-121.95,-19749.,-6281.8,-4216.7,-2607.8,64.119,2284.2,2082.8,1751.3,324.30,3899.9,1686.6,0.0000,7169.2,4449.7,4252.8,3658.0,0.0000,-359.98,-110.95,-92.901,-42.746,-124.98,-587.69,0.0000,-1068.7,-1559.6,-751.83,-1241.6
976.0000000000,89.199,1940.3,2003.3,1699.0,295.73,3701.6,970.66,2.4006,6097.5,2693.3,3357.8,2011.9,0.0000,-6890.9,-6990.4,-1474.2,-2294.8,-2386.4,-16152.,-121.88,-19747.,-6281.4,-4216.1,-2606.9,63.872,2275.4,2074.8,1739.2,322.96,3871.5,1686.6,0.0000,7152.0,4449.7,4252.8,3658.0,0.0000,-358.52,-110.48,-92.364,-42.582,-123.99,-587.69,0.0000,-1068.5,-1559.5,-751.81,-1241.5
977.0000000000,88.965,1933.7,1996.7,1688.2,294.55,3676.6,970.66,2.4012,6082.9,2693.5,3357.9,2012.0,0.0000,-6885.0,-6988.0,-1472.0,-2293.6,-2383.0,-16150.,-121.81,-19745.,-6280.9,-4215.6,-2606.1,63.625,2266.6,2066.8,1727.3,321.62,3843.2,1686.6,0.0000,7134.9,4449.7,4252.8,3658.0,0.0000,-357.05,-110.01,-91.827,-42.417,-123.00,-587.69,0.0000,-1068.4,-1559.4,-751.80,-1241.3
978.0000000000,88.713,1926.7,1989.5,1677.4,293.38,3651.5,970.66,2.4017,6068.0,2693.6,3358.0,2012.1,0.0000,-6878.9,-6985.5,-1469.6,-2292.5,-2379.6,-16148.,-121.74,-19743.,-6280.5,-4215.0,-2605.3,63.374,2257.7,2058.6,1715.3,320.27,3814.9,1686.6,0.0000,7117.7,4449.7,4252.8,3658.0,0.0000,-355.56,-109.53,-91.289,-42.250,-122.01,-587.69,0.0000,-1068.2,-1559.3,-751.78,-1241.2
979.0000000000,88.460,1919.9,1982.3,1666.6,292.20,3626.5,970.49,2.4053,6053.0,2693.7,3358.0,2012.2,0.0000,-6872.6,-6982.9,-1467.2,-2291.3,-2376.0,-16147.,-121.67,-19741.,-6280.0,-4214.4,-2604.5,63.127,2248.9,2050.6,1703.5,318.93,3787.0,1686.6,0.0000,7100.8,4449.7,4252.8,3658.0,0.0000,-354.09,-109.05,-90.757,-42.085,-121.03,-587.69,0.0000,-1068.1,-1559.2,-751.77,-1241.0
980.0000000000,88.208,1913.2,1975.1,1655.7,291.03,3601.8,970.46,2.4122,6037.8,2693.9,3358.0,2012.3,0.0000,-6866.2,-6980.3,-1464.8,-2290.1,-2372.3,-16145.,-121.60,-19739.,-6279.6,-4213.8,-2603.7,62.884,2240.2,2042.7,1691.8,317.61,3759.5,1686.6,0.0000,7084.1,4449.7,4252.8,3658.0,0.0000,-352.64,-108.59,-90.233,-41.923,-120.06,-587.69,0.0000,-1067.9,-1559.1,-751.75,-1240.9
981.0000000000,88.089,1906.2,1968.3,1644.9,289.85,3577.2,970.46,2.5789,6022.6,2694.0,3358.1,2012.5,0.0000,-6859.6,-6977.6,-1462.3,-2288.9,-2368.5,-16143.,-121.53,-19737.,-6279.1,-4213.3,-2602.9,62.641,2231.5,2034.8,1680.2,316.30,3732.1,1686.6,0.0000,7067.5,4449.7,4252.8,3658.0,0.0000,-351.19,-108.12,-89.710,-41.760,-119.09,-587.69,0.0000,-1067.8,-1559.0,-751.74,-1240.8
982.0000000000,87.936,1899.2,1961.8,1634.3,288.69,3552.3,970.46,2.9153,6007.6,2694.1,3358.1,2012.6,0.0000,-6853.0,-6974.9,-1459.8,-2287.7,-2364.7,-16141.,-121.46,-19735.,-6278.6,-4212.7,-2602.1,62.403,2223.1,2027.1,1668.8,315.01,3705.1,1686.6,0.0000,7051.2,4449.7,4252.8,3658.0,0.0000,-349.77,-107.66,-89.198,-41.602,-118.13,-587.69,0.0000,-1067.6,-1558.8,-751.73,-1240.6
983.0000000000,87.921,1892.9,1955.3,1623.8,287.64,3528.2,970.46,2.7944,5992.4,2694.0,3358.2,2012.8,0.0000,-6846.3,-6972.1,-1457.2,-2286.5,-2360.7,-16139.,-121.39,-19733.,-6278.2,-4212.1,-2601.2,62.294,2219.2,2023.5,1666.5,314.42,3694.5,1686.6,2.0606,7045.8,4451.2,4254.2,3658.3,0.0000,-349.07,-107.42,-88.965,-41.530,-117.67,-587.69,-0.94191E-01,-1067.5,-1558.7,-751.72,-1240.5
984.0000000000,87.743,1887.6,1949.7,1614.5,286.79,3506.8,970.45,2.7601,5977.6,2694.0,3358.2,2012.9,0.0000,-6839.7,-6969.4,-1454.7,-2285.3,-2356.8,-16137.,-121.32,-19730.,-6277.7,-4211.5,-2600.4,62.074,2211.4,2016.4,1653.2,313.23,3668.3,1686.6,0.0000,7028.8,4449.7,4252.8,3658.0,0.0000,-347.75,-106.99,-88.494,-41.383,-116.78,-587.69,0.0000,-1067.4,-1558.6,-751.70,-1240.4
985.0000000000,87.553,1882.0,1943.9,1605.7,285.88,3492.3,970.42,2.6006,5963.2,2693.9,3358.3,2013.0,0.0000,-6833.0,-6966.6,-1452.2,-2284.1,-2352.8,-16136.,-121.25,-19728.,-6277.3,-4210.9,-2599.6,61.934,2206.4,2011.8,1645.0,312.45,3648.5,1686.6,0.49303E-01,7016.8,4449.7,4252.8,3658.0,0.0000,-346.87,-106.70,-88.140,-41.289,-116.05,-587.69,-0.22536E-02,-1067.3,-1558.5,-751.68,-1240.2
986.0000000000,87.389,1876.8,1938.8,1597.0,285.11,3470.8,970.42,2.5699,5949.0,2694.0,3358.3,2013.2,0.0000,-6826.4,-6963.8,-1449.7,-2283.0,-2348.8,-16134.,-121.18,-19726.,-6276.8,-4210.4,-2598.8,61.722,2198.8,2005.0,1634.5,311.30,3623.6,1686.6,0.0000,7001.7,4449.7,4252.8,3658.0,0.0000,-345.60,-106.29,-87.673,-41.148,-115.16,-587.69,0.0000,-1067.1,-1558.4,-751.67,-1240.1
987.0000000000,87.205,1871.0,1933.1,1588.2,284.16,3449.1,970.42,2.5704,5934.8,2694.1,3358.4,2013.3,0.0000,-6819.7,-6961.0,-1447.1,-2281.8,-2344.8,-16132.,-121.11,-19724.,-6276.3,-4209.8,-2598.0,61.517,2191.5,1998.3,1624.2,310.18,3599.1,1686.6,0.0000,6986.9,4449.7,4252.8,3658.0,0.0000,-344.36,-105.88,-87.213,-41.011,-114.28,-587.69,0.0000,-1067.0,-1558.3,-751.65,-1239.9
988.0000000000,86.999,1864.8,1927.0,1579.1,283.23,3427.2,970.42,2.4203,5921.0,2694.2,3358.4,2013.4,0.0000,-6813.0,-6958.1,-1444.6,-2280.6,-2340.6,-16130.,-121.04,-19721.,-6275.9,-4209.2,-2597.2,61.314,2184.3,1991.7,1613.9,309.07,3574.8,1686.6,0.0000,6972.1,4449.7,4252.8,3658.0,0.0000,-343.13,-105.48,-86.758,-40.876,-113.40,-587.69,0.0000,-1066.8,-1558.2,-751.64,-1239.8
989.0000000000,86.803,1859.0,1920.8,1569.8,282.26,3405.2,970.42,2.4065,5907.7,2694.3,3358.4,2013.7,0.0000,-6806.2,-6955.3,-1442.0,-2279.4,-2336.4,-16128.,-120.97,-19719.,-6275.4,-4208.6,-2596.4,61.110,2177.0,1985.1,1603.7,307.96,3550.5,1686.6,0.0000,6957.4,4449.7,4252.8,3658.0,0.0000,-341.90,-105.08,-86.303,-40.740,-112.52,-587.69,0.0000,-1066.7,-1558.1,-751.62,-1239.7
990.0000000000,86.593,1853.1,1914.9,1560.2,281.29,3384.1,970.42,2.4070,5895.3,2694.4,3358.4,2013.8,0.0000,-6799.4,-6952.5,-1439.4,-2278.1,-2332.1,-16126.,-120.90,-19717.,-6274.9,-4208.0,-2595.6,60.907,2169.8,1978.5,1593.5,306.85,3526.3,1686.6,0.0000,6942.7,4449.7,4252.8,3658.0,0.0000,-340.67,-104.68,-85.850,-40.605,-111.65,-587.69,0.0000,-1066.5,-1558.0,-751.61,-1239.5
991.0000000000,86.385,1847.0,1909.0,1550.5,280.31,3363.1,970.42,2.4076,5882.6,2694.5,3358.4,2014.0,0.0000,-6792.5,-6949.7,-1436.8,-2276.9,-2327.7,-16124.,-120.83,-19714.,-6274.5,-4207.4,-2594.8,60.701,2162.4,1971.8,1583.3,305.73,3502.1,1686.6,0.0000,6928.1,4449.7,4252.8,3658.0,0.0000,-339.43,-104.28,-85.395,-40.467,-110.77,-587.69,0.0000,-1066.4,-1557.9,-751.59,-1239.4
992.0000000000,86.176,1841.0,1902.7,1540.9,279.34,3341.9,970.41,2.3537,5869.7,2694.6,3358.4,2014.1,0.0000,-6785.6,-6946.8,-1434.1,-2275.7,-2323.2,-16122.,-120.76,-19712.,-6274.0,-4206.9,-2593.9,60.497,2155.2,1965.2,1573.2,304.63,3478.2,1686.6,0.0000,6913.6,4449.7,4252.8,3658.0,0.0000,-338.19,-103.88,-84.944,-40.331,-109.90,-587.69,0.0000,-1066.2,-1557.8,-751.58,-1239.2
993.0000000000,85.968,1835.0,1896.6,1531.5,278.38,3320.4,970.38,2.2174,5856.4,2694.7,3358.5,2014.2,0.0000,-6778.6,-6944.0,-1431.4,-2274.5,-2318.7,-16120.,-120.69,-19710.,-6273.6,-4206.3,-2593.1,60.301,2148.2,1958.8,1563.4,303.56,3454.8,1686.6,0.0000,6899.4,4449.7,4252.8,3658.0,0.0000,-337.01,-103.49,-84.506,-40.201,-109.05,-587.69,0.0000,-1066.1,-1557.7,-751.57,-1239.1
994.0000000000,85.764,1829.2,1890.4,1522.0,277.44,3298.6,970.38,2.2179,5842.8,2694.8,3358.5,2014.3,0.0000,-6771.5,-6941.1,-1428.7,-2273.3,-2314.2,-16118.,-120.63,-19707.,-6273.1,-4205.7,-2592.3,60.112,2141.4,1952.6,1553.7,302.52,3431.7,1686.6,0.0000,6885.4,4449.7,4252.8,3658.0,0.0000,-335.85,-103.11,-84.077,-40.074,-108.20,-587.69,0.0000,-1065.9,-1557.6,-751.55,-1239.0
995.0000000000,85.563,1823.5,1884.0,1512.7,276.51,3277.0,970.38,2.2184,5829.4,2694.9,3358.5,2014.5,0.0000,-6764.5,-6938.2,-1426.0,-2272.0,-2309.5,-16116.,-120.56,-19705.,-6272.6,-4205.1,-2591.5,59.925,2134.8,1946.6,1544.1,301.50,3409.0,1686.6,0.0000,6871.6,4449.7,4252.8,3658.0,0.0000,-334.72,-102.74,-83.654,-39.950,-107.37,-587.69,0.0000,-1065.8,-1557.5,-751.54,-1238.8
996.0000000000,85.367,1817.9,1878.2,1503.5,275.52,3255.7,970.38,2.2189,5816.1,2695.0,3358.5,2014.6,0.0000,-6757.4,-6935.4,-1423.2,-2270.8,-2304.9,-16114.,-120.49,-19702.,-6272.2,-4204.5,-2590.7,59.744,2128.3,1940.7,1534.7,300.51,3386.6,1686.6,0.0000,6858.0,4449.7,4252.8,3658.0,0.0000,-333.61,-102.38,-83.239,-39.829,-106.55,-587.69,0.0000,-1065.6,-1557.4,-751.52,-1238.7
997.0000000000,85.176,1812.5,1872.7,1494.4,274.61,3234.8,970.37,2.2194,5802.8,2695.0,3358.6,2014.7,0.0000,-6750.3,-6932.5,-1420.5,-2269.6,-2300.2,-16112.,-120.42,-19700.,-6271.7,-4203.9,-2589.9,59.572,2122.2,1935.1,1525.6,299.57,3364.9,1686.6,0.0000,6844.8,4449.7,4252.8,3658.0,0.0000,-332.55,-102.04,-82.838,-39.715,-105.75,-587.69,0.0000,-1065.5,-1557.3,-751.51,-1238.6
998.0000000000,85.080,1807.4,1867.2,1485.4,273.76,3214.0,970.37,2.0808,5789.6,2695.0,3358.6,2014.9,0.0000,-6743.2,-6929.7,-1417.7,-2268.4,-2295.5,-16110.,-120.35,-19697.,-6271.3,-4203.3,-2589.1,59.407,2116.3,1929.8,1516.6,298.65,3343.5,1686.6,0.0000,6831.9,4449.7,4252.8,3658.0,0.0000,-331.54,-101.70,-82.447,-39.605,-104.96,-587.69,0.0000,-1065.4,-1557.2,-751.49,-1238.4
999.0000000000,84.814,1802.2,1861.8,1476.5,272.94,3193.4,970.33,2.0513,5776.6,2695.1,3358.6,2015.0,0.0000,-6736.1,-6926.8,-1414.9,-2267.1,-2290.7,-16108.,-120.28,-19695.,-6270.8,-4202.7,-2588.3,59.246,2110.6,1924.5,1507.8,297.77,3322.5,1686.6,0.0000,6819.1,4449.7,4252.8,3658.0,0.0000,-330.55,-101.38,-82.063,-39.497,-104.18,-587.69,0.0000,-1065.2,-1557.1,-751.48,-1238.3
1000.000000000,84.642,1797.5,1856.6,1467.9,272.20,3173.2,970.33,2.0518,5763.7,2695.2,3358.6,2015.1,0.0000,-6729.0,-6924.0,-1412.1,-2265.9,-2286.0,-16106.,-120.21,-19692.,-6270.3,-4202.1,-2587.5,59.177,2108.2,1922.3,1501.3,297.34,3306.3,1686.6,0.0000,6809.3,4449.7,4252.8,3658.0,0.0000,-330.07,-101.21,-81.804,-39.452,-103.55,-587.69,0.0000,-1065.1,-1556.9,-751.46,-1238.1
1001.000000000,84.517,1793.7,1852.3,1459.6,271.59,3153.9,970.31,2.0523,5751.1,2695.1,3358.5,2015.2,0.0000,-6722.0,-6921.3,-1409.4,-2264.7,-2281.2,-16104.,-120.15,-19690.,-6269.9,-4201.5,-2586.7,59.022,2102.6,1917.2,1492.7,296.48,3285.8,1686.6,0.0000,6796.8,4449.7,4252.8,3658.0,0.0000,-329.11,-100.89,-81.431,-39.348,-102.79,-587.69,0.0000,-1065.0,-1556.8,-751.45,-1238.0
1002.000000000,84.372,1789.5,1847.8,1451.6,270.86,3134.8,970.29,2.0528,5738.9,2695.2,3358.5,2015.4,0.0000,-6715.0,-6918.6,-1406.6,-2263.5,-2276.4,-16102.,-120.08,-19687.,-6269.4,-4200.9,-2585.9,58.868,2097.1,1912.2,1484.2,295.63,3265.4,1686.6,0.0000,6784.5,4449.7,4252.8,3658.0,0.0000,-328.16,-100.58,-81.061,-39.245,-102.03,-587.69,0.0000,-1064.8,-1556.7,-751.43,-1237.9
1003.000000000,84.219,1785.0,1842.9,1443.6,270.19,3115.8,970.29,2.0533,5726.8,2695.3,3358.5,2015.5,0.0000,-6708.0,-6915.9,-1403.9,-2262.3,-2271.6,-16100.,-120.01,-19685.,-6269.0,-4200.4,-2585.1,58.716,2091.7,1907.3,1475.8,294.78,3245.3,1686.6,0.0000,6772.3,4449.7,4252.8,3658.0,0.0000,-327.22,-100.27,-80.695,-39.144,-101.27,-587.69,0.0000,-1064.7,-1556.6,-751.42,-1237.7
1004.000000000,83.916,1780.6,1838.3,1435.6,269.45,3096.8,970.29,2.0538,5714.7,2695.3,3358.5,2015.6,0.0000,-6701.0,-6913.3,-1401.1,-2261.1,-2266.8,-16098.,-119.94,-19682.,-6268.5,-4199.8,-2584.3,58.549,2085.8,1901.9,1467.1,293.87,3224.6,1686.6,0.0000,6759.7,4449.7,4252.8,3658.0,0.0000,-326.19,-99.938,-80.311,-39.033,-100.50,-587.69,0.0000,-1064.6,-1556.5,-751.40,-1237.6
1005.000000000,83.644,1776.1,1833.4,1427.5,268.67,3077.7,970.27,2.0549,5703.0,2695.4,3358.5,2015.8,0.0000,-6694.1,-6910.7,-1398.3,-2259.9,-2261.9,-16096.,-119.88,-19680.,-6268.1,-4199.2,-2583.5,58.380,2079.8,1896.4,1458.5,292.94,3203.9,1686.6,0.0000,6747.2,4449.7,4252.8,3658.0,0.0000,-325.16,-99.601,-79.927,-38.920,-99.734,-587.69,0.0000,-1064.4,-1556.4,-751.39,-1237.5
1006.000000000,83.476,1771.3,1828.3,1419.5,267.89,3058.8,970.25,2.0599,5691.3,2695.5,3358.6,2015.9,0.0000,-6687.1,-6908.0,-1395.5,-2258.7,-2257.1,-16094.,-119.81,-19677.,-6267.6,-4198.6,-2582.7,58.222,2074.1,1891.2,1450.1,292.07,3183.9,1686.6,0.0000,6735.1,4449.7,4252.8,3658.0,0.0000,-324.18,-99.282,-79.558,-38.814,-98.984,-587.69,0.0000,-1064.3,-1556.3,-751.37,-1237.3
1007.000000000,83.321,1766.6,1823.4,1411.4,267.11,3040.1,970.25,2.0603,5680.0,2695.6,3358.6,2016.0,0.0000,-6680.1,-6905.3,-1392.7,-2257.5,-2252.2,-16092.,-119.74,-19675.,-6267.1,-4198.0,-2581.9,58.070,2068.7,1886.3,1441.9,291.24,3164.3,1686.6,0.0000,6723.2,4449.7,4252.8,3658.0,0.0000,-323.25,-98.975,-79.199,-38.713,-98.248,-587.69,0.0000,-1064.2,-1556.2,-751.36,-1237.2
1008.000000000,83.040,1762.2,1818.5,1403.3,266.36,3021.8,970.25,2.0608,5668.6,2695.7,3358.6,2016.1,0.0000,-6673.1,-6902.6,-1389.9,-2256.3,-2247.3,-16090.,-119.67,-19672.,-6266.7,-4197.4,-2581.1,57.924,2063.5,1881.6,1433.8,290.43,3145.1,1686.6,0.0000,6711.5,4449.7,4252.8,3658.0,0.0000,-322.34,-98.679,-78.849,-38.616,-97.525,-587.69,0.0000,-1064.0,-1556.1,-751.34,-1237.0
1009.000000000,82.882,1758.0,1813.7,1395.3,265.64,3003.7,970.25,2.0613,5657.3,2695.9,3358.6,2016.2,0.0000,-6666.2,-6900.0,-1387.1,-2255.0,-2242.4,-16088.,-119.61,-19670.,-6266.2,-4196.8,-2580.3,57.787,2058.6,1877.1,1426.0,289.67,3126.4,1686.6,0.0000,6700.2,4449.7,4252.8,3658.0,0.0000,-321.49,-98.398,-78.512,-38.525,-96.817,-587.69,0.0000,-1063.9,-1556.0,-751.33,-1236.9
1010.000000000,82.732,1753.9,1809.2,1387.6,264.94,2985.6,970.25,1.9952,5645.9,2696.0,3358.6,2016.4,0.0000,-6659.3,-6897.4,-1384.3,-2253.8,-2237.6,-16086.,-119.54,-19667.,-6265.8,-4196.1,-2579.5,57.645,2053.6,1872.5,1418.2,288.88,3107.6,1686.6,0.0000,6688.8,4449.7,4252.8,3658.0,0.0000,-320.61,-98.109,-78.170,-38.430,-96.107,-587.69,0.0000,-1063.8,-1555.9,-751.31,-1236.8
1011.000000000,82.573,1749.8,1804.5,1379.9,264.25,2967.6,970.25,1.8783,5634.7,2696.1,3358.6,2016.5,0.0000,-6652.4,-6894.7,-1381.5,-2252.6,-2232.7,-16084.,-119.48,-19664.,-6265.3,-4195.5,-2578.7,57.503,2048.5,1867.9,1410.4,288.09,3088.8,1686.6,0.0000,6677.4,4449.7,4252.8,3658.0,0.0000,-319.72,-97.819,-77.829,-38.335,-95.399,-587.69,0.0000,-1063.6,-1555.8,-751.30,-1236.6
1012.000000000,82.492,1747.8,1801.8,1372.7,263.90,2951.2,970.23,1.8872,5623.5,2696.2,3358.6,2016.7,0.0000,-6645.7,-6892.2,-1378.8,-2251.4,-2227.9,-16082.,-119.41,-19662.,-6264.9,-4194.9,-2577.9,57.986,2062.2,1880.6,1423.0,290.35,3115.5,1686.6,4.0531,6694.0,4450.6,4253.7,3658.5,0.0000,-321.69,-98.417,-78.413,-38.583,-96.109,-587.69,-0.18523,-1063.7,-1555.7,-751.29,-1236.5
1013.000000000,82.689,1750.5,1803.7,1368.0,264.33,2939.4,970.23,1.8877,5613.7,2696.3,3358.6,2016.8,0.0000,-6639.5,-6890.0,-1376.2,-2250.3,-2223.3,-16080.,-119.35,-19659.,-6264.4,-4194.3,-2577.1,58.042,2073.7,1885.4,1431.3,290.74,3113.7,1686.6,107.35,6699.0,4458.2,4262.5,3673.9,0.0000,-322.56,-98.651,-78.449,-38.695,-95.830,-587.69,-4.9059,-1063.8,-1555.6,-751.32,-1236.8
1014.000000000,82.795,1753.5,1805.7,1365.7,264.69,2930.1,970.22,1.8882,5605.0,2696.5,3358.6,2016.9,0.0000,-6633.7,-6888.1,-1373.7,-2249.2,-2218.9,-16077.,-119.29,-19657.,-6264.0,-4193.7,-2576.3,58.036,2067.5,1885.2,1414.7,290.61,3094.6,1686.6,0.0000,6680.8,4457.2,4262.6,3673.0,0.0000,-322.43,-98.602,-78.252,-38.690,-95.233,-587.69,0.0000,-1063.5,-1555.5,-751.30,-1236.6
1015.000000000,82.807,1754.3,1805.8,1362.7,264.89,2919.4,970.19,1.8887,5596.6,2696.6,3358.6,2017.0,0.0000,-6628.2,-6886.2,-1371.3,-2248.2,-2214.7,-16075.,-119.23,-19654.,-6263.5,-4193.1,-2575.5,57.954,2064.6,1882.5,1407.6,290.12,3076.8,1686.6,0.0000,6670.0,4453.5,4257.3,3664.6,0.0000,-321.90,-98.424,-77.966,-38.636,-94.565,-587.69,0.0000,-1063.4,-1555.4,-751.26,-1236.3
1016.000000000,82.876,1753.0,1804.5,1359.7,264.75,2906.9,970.19,1.8892,5587.7,2696.7,3358.6,2017.1,0.0000,-6622.7,-6884.3,-1368.8,-2247.1,-2210.5,-16073.,-119.17,-19652.,-6263.1,-4192.5,-2574.7,57.844,2060.7,1879.0,1400.2,289.49,3058.7,1686.6,0.0000,6659.0,4451.0,4254.4,3660.2,0.0000,-321.21,-98.200,-77.656,-38.563,-93.885,-587.69,0.0000,-1063.3,-1555.3,-751.23,-1236.0
1017.000000000,82.850,1750.5,1802.4,1354.8,264.33,2893.3,970.19,1.8898,5578.8,2696.8,3358.6,2017.3,0.0000,-6617.1,-6882.4,-1366.4,-2246.0,-2206.3,-16071.,-119.11,-19649.,-6262.6,-4191.9,-2573.9,57.735,2056.8,1875.4,1393.0,288.86,3041.1,1686.6,0.0000,6648.3,4450.1,4253.3,3658.6,0.0000,-320.52,-97.976,-77.352,-38.490,-93.221,-587.69,0.0000,-1063.1,-1555.2,-751.21,-1235.8
1018.000000000,82.765,1747.8,1799.7,1349.5,263.82,2878.5,970.19,1.8932,5570.4,2696.9,3358.6,2017.4,0.0000,-6611.6,-6880.5,-1364.0,-2244.9,-2202.2,-16069.,-119.05,-19647.,-6262.2,-4191.3,-2573.1,57.616,2052.5,1871.6,1385.7,288.19,3023.5,1686.6,0.0000,6637.6,4449.8,4252.9,3658.1,0.0000,-319.79,-97.737,-77.043,-38.411,-92.556,-587.69,0.0000,-1063.0,-1555.1,-751.19,-1235.7
1019.000000000,82.694,1744.9,1797.1,1343.3,263.26,2864.2,970.17,1.8937,5563.7,2697.0,3358.6,2017.5,0.0000,-6605.9,-6878.5,-1361.5,-2243.8,-2198.1,-16067.,-118.99,-19644.,-6261.7,-4190.7,-2572.3,57.500,2048.4,1867.8,1378.6,287.53,3006.3,1686.6,0.0000,6627.2,4449.7,4252.8,3658.0,0.0000,-319.06,-97.502,-76.739,-38.333,-91.903,-587.69,0.0000,-1062.9,-1555.0,-751.17,-1235.6
1020.000000000,82.707,1741.5,1794.2,1336.6,262.66,2852.0,970.17,1.8942,5558.3,2697.1,3358.7,2017.6,0.0000,-6600.3,-6876.5,-1359.0,-2242.7,-2194.1,-16065.,-118.93,-19641.,-6261.3,-4190.1,-2571.5,57.389,2044.5,1864.2,1371.7,286.91,2989.6,1686.6,0.0000,6617.1,4449.7,4252.8,3658.0,0.0000,-318.37,-97.277,-76.445,-38.260,-91.265,-587.69,0.0000,-1062.7,-1554.9,-751.16,-1235.4
1021.000000000,82.590,1738.7,1791.4,1329.7,262.00,2840.5,970.17,1.8947,5551.7,2697.2,3358.7,2017.8,0.0000,-6594.7,-6874.5,-1356.5,-2241.6,-2190.2,-16063.,-118.87,-19639.,-6260.8,-4189.5,-2570.7,57.282,2040.6,1860.7,1364.9,286.30,2973.2,1686.6,0.0000,6607.1,4449.7,4252.8,3658.0,0.0000,-317.70,-97.057,-76.158,-38.188,-90.638,-587.69,0.0000,-1062.6,-1554.8,-751.14,-1235.3
1022.000000000,82.474,1735.9,1788.3,1323.4,261.45,2827.5,970.17,1.8702,5543.9,2697.3,3358.7,2017.9,0.0000,-6589.1,-6872.5,-1353.9,-2240.5,-2186.4,-16060.,-118.81,-19636.,-6260.4,-4188.8,-2569.9,57.175,2036.8,1857.2,1358.2,285.69,2957.0,1686.6,0.0000,6597.3,4449.7,4252.8,3658.0,0.0000,-317.03,-96.839,-75.874,-38.117,-90.017,-587.69,0.0000,-1062.5,-1554.7,-751.13,-1235.2
1023.000000000,82.360,1732.8,1785.0,1317.4,260.91,2812.9,970.17,1.7258,5535.1,2697.5,3358.8,2018.1,0.0000,-6583.5,-6870.5,-1351.3,-2239.4,-2182.6,-16058.,-118.75,-19634.,-6259.9,-4188.2,-2569.1,57.069,2033.1,1853.8,1351.6,285.10,2941.0,1686.6,0.0000,6587.6,4449.7,4252.8,3658.0,0.0000,-316.37,-96.621,-75.593,-38.046,-89.393,-587.69,0.0000,-1062.4,-1554.6,-751.11,-1235.0
1024.000000000,82.248,1729.8,1781.8,1311.2,260.37,2797.6,970.17,1.7263,5525.8,2697.6,3358.8,2018.2,0.0000,-6577.8,-6868.5,-1348.7,-2238.3,-2178.8,-16056.,-118.69,-19631.,-6259.5,-4187.6,-2568.3,56.961,2029.2,1850.3,1344.9,284.48,2925.0,1686.6,0.0000,6577.9,4449.7,4252.8,3658.0,0.0000,-315.69,-96.400,-75.311,-37.974,-88.764,-587.69,0.0000,-1062.3,-1554.5,-751.10,-1234.9
1025.000000000,82.088,1727.1,1778.7,1304.8,259.86,2782.4,970.17,1.7268,5516.1,2697.7,3358.8,2018.3,0.0000,-6572.2,-6866.5,-1346.1,-2237.1,-2174.9,-16054.,-118.63,-19629.,-6259.0,-4187.0,-2567.5,56.892,2026.7,1848.1,1339.6,284.08,2912.0,1686.6,0.0000,6570.0,4449.7,4252.8,3658.0,0.0000,-315.23,-96.247,-75.093,-37.928,-88.225,-587.69,0.0000,-1062.2,-1554.4,-751.08,-1234.8
1026.000000000,81.732,1725.6,1776.9,1298.6,259.59,2768.0,970.15,1.7272,5506.6,2697.8,3358.8,2018.5,0.0000,-6566.7,-6864.6,-1343.5,-2236.1,-2171.1,-16052.,-118.58,-19626.,-6258.6,-4186.4,-2566.7,57.301,2033.9,1855.4,1335.9,284.84,2900.2,1686.6,0.0000,6562.8,4449.7,4252.8,3658.0,0.0000,-316.15,-96.546,-75.056,-38.047,-87.723,-587.69,0.0000,-1062.0,-1554.3,-751.07,-1234.6
1027.000000000,81.648,1746.3,1795.2,1293.8,262.95,2757.8,970.13,1.7324,5498.2,2697.9,3358.8,2018.6,0.0000,-6563.0,-6863.8,-1341.2,-2235.1,-2167.3,-16049.,-118.52,-19623.,-6258.1,-4185.8,-2565.9,79.639,2245.1,2071.9,1401.8,311.27,3005.5,1687.0,436.32,6629.5,4461.9,4267.1,3679.9,0.0000,-342.37,-105.88,-79.507,-41.224,-90.692,-587.69,-19.938,-1062.5,-1554.2,-751.12,-1235.1
1028.000000000,83.887,1813.8,1853.4,1317.1,274.06,2824.4,970.13,1.7350,5503.3,2698.0,3358.8,2018.7,0.0000,-6564.5,-6865.8,-1342.1,-2234.8,-2165.7,-16047.,-118.47,-19621.,-6257.7,-4185.1,-2565.2,890.83,3461.4,3000.6,2058.0,384.87,4639.2,1701.6,1043.1,7631.2,4531.8,4380.3,3873.9,0.0000,-361.43,-128.84,-102.61,-43.603,-140.59,-587.92,-47.664,-1069.7,-1554.1,-751.69,-1239.9
1029.000000000,86.415,1886.8,1923.6,1448.3,286.66,3066.9,970.13,1.7355,5559.1,2698.1,3358.8,2018.9,0.0000,-6570.3,-6870.4,-1347.4,-2235.0,-2169.1,-16045.,-118.42,-19619.,-6257.3,-4184.5,-2564.4,66.665,2374.9,2165.5,2079.4,530.93,4666.7,1686.7,0.0000,7700.2,4497.7,4416.6,3797.9,0.0000,-369.28,-112.82,-103.77,-45.616,-140.78,-587.69,0.0000,-1070.7,-1554.0,-751.87,-1237.9
1030.000000000,88.281,1937.2,1974.5,1606.8,302.77,3317.3,970.09,1.7360,5639.1,2698.0,3359.2,2019.0,0.0000,-6578.1,-6876.0,-1354.4,-2235.2,-2178.5,-16043.,-118.37,-19618.,-6256.8,-4183.9,-2563.6,66.976,2386.0,2175.6,2046.7,369.75,4618.0,1686.6,0.0000,7607.4,4480.8,4289.6,3695.4,0.0000,-371.05,-113.41,-103.98,-44.821,-140.65,-587.69,0.0000,-1069.3,-1553.9,-751.19,-1235.1
1031.000000000,90.257,1962.6,2002.5,1722.1,308.18,3460.6,970.04,1.7365,5698.0,2698.1,3359.0,2019.5,0.0000,-6586.3,-6881.2,-1362.4,-2235.4,-2187.4,-16041.,-118.31,-19617.,-6256.4,-4183.3,-2562.8,67.037,2388.2,2177.6,2038.9,356.62,4606.7,1686.6,0.0000,7599.3,4464.4,4271.4,3676.8,0.0000,-371.45,-113.58,-104.02,-44.778,-140.76,-587.69,0.0000,-1069.2,-1553.8,-751.09,-1234.5
1032.000000000,90.730,1974.6,2019.1,1802.9,310.52,3558.2,970.04,1.7370,5740.0,2698.2,3359.1,2019.8,0.0000,-6593.8,-6885.7,-1370.2,-2235.4,-2193.6,-16039.,-118.25,-19616.,-6255.9,-4182.7,-2562.0,67.001,2386.9,2176.4,2034.8,348.23,4600.8,1686.6,0.0000,7594.8,4456.1,4260.8,3666.0,0.0000,-371.31,-113.58,-103.99,-44.704,-140.91,-587.69,0.0000,-1069.1,-1553.7,-751.01,-1234.1
1033.000000000,91.051,1982.4,2027.2,1853.1,310.99,3614.4,970.05,1.7375,5811.4,2698.3,3359.3,2020.2,0.0000,-6600.3,-6889.6,-1380.7,-2235.3,-2198.4,-16037.,-118.20,-19614.,-6255.5,-4182.0,-2561.2,67.045,2388.4,2177.9,2033.1,344.59,4598.0,1686.6,0.0000,7593.0,4451.9,4255.6,3660.7,0.0000,-371.62,-113.72,-104.02,-44.709,-141.06,-587.69,0.0000,-1069.1,-1553.6,-750.97,-1233.8
1034.000000000,91.139,1995.4,2041.3,1873.9,312.37,3679.8,970.05,1.6077,5932.2,2698.4,3359.3,2020.3,0.0000,-6606.8,-6893.4,-1388.1,-2235.1,-2202.2,-16035.,-118.14,-19614.,-6255.1,-4181.4,-2560.4,821.51,3472.9,2600.4,2159.3,516.12,4741.9,1686.6,2397.6,7738.4,4613.7,4448.9,3872.3,0.0000,-381.66,-124.30,-105.02,-46.721,-141.90,-587.69,-109.56,-1071.2,-1553.5,-751.96,-1239.1
1035.000000000,91.940,2019.7,2067.8,1877.6,315.62,3838.6,970.05,1.5688,6098.8,2698.5,3359.5,2020.7,0.0000,-6614.3,-6897.7,-1393.7,-2235.1,-2205.5,-16033.,-118.09,-19613.,-6254.6,-4180.8,-2559.7,69.141,2463.1,2245.9,2136.7,353.34,4616.9,1686.6,0.0000,7823.5,4744.9,4368.8,3845.0,0.0000,-383.42,-117.42,-105.42,-46.100,-141.45,-587.69,0.0000,-1072.4,-1553.4,-751.53,-1238.3
1036.000000000,92.455,2042.6,2091.8,1879.9,317.40,3991.3,970.05,29.355,6191.9,2698.6,3360.0,2022.2,0.0000,-6622.6,-6902.2,-1398.3,-2235.1,-2208.3,-16031.,-118.03,-19613.,-6254.2,-4180.2,-2558.9,69.228,2466.2,2248.8,2071.7,353.35,4601.9,1686.6,0.0000,7662.3,4557.0,4270.3,3680.4,0.0000,-383.99,-117.64,-105.48,-46.156,-141.49,-587.69,0.0000,-1070.1,-1553.3,-751.00,-1233.9
1037.000000000,92.875,2053.1,2102.4,1901.4,319.17,4040.6,970.05,46.226,6241.1,2699.0,3361.0,2024.9,0.0000,-6630.6,-6906.3,-1402.3,-2235.0,-2210.9,-16029.,-117.98,-19612.,-6253.7,-4179.6,-2558.1,69.179,2464.4,2247.2,2055.9,352.57,4598.8,1686.6,0.0000,7627.3,4501.5,4260.7,3668.8,0.0000,-383.81,-117.63,-105.45,-46.119,-141.58,-587.69,0.0000,-1069.6,-1553.2,-750.94,-1233.5
1038.000000000,92.797,2056.8,2106.0,1917.5,319.68,4054.3,970.05,50.844,6260.5,2701.7,3362.0,2024.4,0.0000,-6637.6,-6910.0,-1405.8,-2234.9,-2213.5,-16027.,-117.93,-19612.,-6253.3,-4179.0,-2557.3,69.063,2460.3,2243.4,2047.3,351.96,4597.6,1686.6,0.0000,7608.5,4474.1,4255.4,3661.8,0.0000,-383.26,-117.50,-105.37,-46.042,-141.67,-587.69,0.0000,-1069.3,-1553.1,-750.89,-1233.2
1039.000000000,92.777,2061.4,2107.3,1920.7,319.43,4052.5,970.05,36.797,6261.9,2702.7,3363.6,2023.9,0.0000,-6643.7,-6913.2,-1409.0,-2234.7,-2216.1,-16025.,-117.87,-19612.,-6252.9,-4178.4,-2556.5,68.907,2454.8,2238.4,2042.4,351.23,4597.2,1686.6,0.0000,7598.9,4460.3,4253.2,3658.8,0.0000,-382.48,-117.29,-105.26,-45.938,-141.76,-587.69,0.0000,-1069.2,-1553.0,-750.87,-1233.0
1040.000000000,92.673,2062.8,2109.4,1920.8,318.91,4066.9,970.06,47.849,6262.3,2703.1,3362.5,2023.5,0.0000,-6648.8,-6916.1,-1411.9,-2234.5,-2218.9,-16023.,-117.82,-19612.,-6252.5,-4177.8,-2555.8,68.738,2448.7,2232.8,2040.1,350.44,4597.2,1686.6,0.0000,7594.2,4453.4,4252.8,3658.0,0.0000,-381.61,-117.06,-105.15,-45.825,-141.85,-587.69,0.0000,-1069.1,-1552.9,-750.85,-1232.9
1041.000000000,92.526,2060.3,2110.0,1920.2,318.27,4090.5,970.05,40.879,6281.7,2704.0,3361.6,2023.9,0.0000,-6653.3,-6918.7,-1414.5,-2234.2,-2222.1,-16022.,-117.76,-19612.,-6252.1,-4177.2,-2555.0,68.628,2444.8,2229.3,2039.2,349.93,4597.1,1686.6,0.0000,7592.6,4450.5,4252.8,3658.0,0.0000,-381.07,-116.92,-105.08,-45.752,-141.94,-587.69,0.0000,-1069.1,-1552.8,-750.84,-1232.7
1042.000000000,92.517,2060.2,2110.4,1925.1,317.74,4121.8,970.03,35.358,6291.4,2706.5,3361.2,2023.4,0.0000,-6657.5,-6921.1,-1417.0,-2233.9,-2225.6,-16020.,-117.71,-19612.,-6251.8,-4176.6,-2554.2,68.495,2440.1,2225.0,2038.6,349.30,4597.1,1686.6,0.0000,7592.4,4450.0,4252.8,3658.0,0.0000,-380.40,-116.73,-104.99,-45.663,-142.02,-587.69,0.0000,-1069.1,-1552.7,-750.83,-1232.6
1043.000000000,92.432,2057.9,2112.5,1930.9,317.15,4130.0,970.03,35.354,6290.2,2705.5,3361.6,2023.2,0.0000,-6661.5,-6923.2,-1419.2,-2233.5,-2229.1,-16018.,-117.65,-19612.,-6251.5,-4176.0,-2553.5,68.321,2433.9,2219.3,2037.8,348.50,4597.0,1686.6,0.0000,7592.3,4450.0,4252.8,3658.0,0.0000,-379.49,-116.48,-104.87,-45.547,-142.10,-587.69,0.0000,-1069.1,-1552.6,-750.81,-1232.5
1044.000000000,92.273,2055.4,2109.2,1930.9,316.52,4132.6,970.03,42.100,6296.6,2704.7,3361.4,2023.2,0.0000,-6665.0,-6925.0,-1421.3,-2233.1,-2232.6,-16016.,-117.59,-19612.,-6251.2,-4175.4,-2552.7,68.136,2427.3,2213.3,2037.0,347.63,4596.9,1686.6,0.0000,7592.3,4449.7,4252.8,3658.0,0.0000,-378.52,-116.20,-104.75,-45.424,-142.18,-587.69,0.0000,-1069.1,-1552.5,-750.80,-1232.4
1045.000000000,92.105,2053.7,2104.9,1930.3,315.90,4131.4,970.04,41.372,6310.0,2704.2,3360.9,2023.3,0.0000,-6667.8,-6926.5,-1423.2,-2232.7,-2236.0,-16015.,-117.54,-19612.,-6250.9,-4174.8,-2551.9,67.945,2420.5,2207.1,2036.1,346.74,4596.8,1686.6,0.0000,7592.3,4449.7,4252.8,3658.0,0.0000,-377.51,-115.90,-104.62,-45.297,-142.25,-587.69,0.0000,-1069.1,-1552.5,-750.79,-1232.2
1046.000000000,91.921,2049.5,2100.6,1929.6,315.20,4144.2,970.04,35.984,6315.3,2703.6,3360.6,2023.3,0.0000,-6670.1,-6927.7,-1424.9,-2232.3,-2239.7,-16013.,-117.48,-19612.,-6250.6,-4174.3,-2551.2,67.761,2414.0,2201.1,2035.3,345.88,4596.8,1686.6,0.0000,7592.2,4449.7,4252.8,3658.0,0.0000,-376.53,-115.61,-104.50,-45.174,-142.33,-587.69,0.0000,-1069.1,-1552.4,-750.77,-1232.1
1047.000000000,91.737,2044.6,2095.6,1929.5,314.59,4145.0,970.02,34.800,6320.1,2703.1,3360.6,2023.2,0.0000,-6671.9,-6928.7,-1426.6,-2231.8,-2243.5,-16011.,-117.43,-19612.,-6250.2,-4173.7,-2550.4,67.586,2407.7,2195.4,2034.5,345.07,4596.7,1686.6,0.0000,7592.2,4449.7,4252.8,3658.0,0.0000,-375.59,-115.33,-104.38,-45.058,-142.40,-587.69,0.0000,-1069.1,-1552.3,-750.76,-1232.0
1048.000000000,91.752,2040.1,2091.4,1929.6,313.86,4153.4,969.99,28.331,6323.7,2702.8,3360.5,2023.2,0.0000,-6673.4,-6929.5,-1428.1,-2231.3,-2247.1,-16010.,-117.37,-19612.,-6249.9,-4173.1,-2549.6,67.454,2403.0,2191.1,2033.9,344.45,4596.6,1686.6,0.0000,7592.2,4449.7,4252.8,3658.0,0.0000,-374.89,-115.13,-104.29,-44.969,-142.47,-587.69,0.0000,-1069.1,-1552.2,-750.75,-1231.8
1049.000000000,91.592,2037.1,2087.5,1928.9,313.30,4164.6,969.99,28.328,6336.3,2702.4,3360.3,2023.2,0.0000,-6674.6,-6930.1,-1429.5,-2230.8,-2250.5,-16008.,-117.32,-19611.,-6249.5,-4172.5,-2548.9,67.399,2401.0,2189.4,2033.6,344.19,4596.6,1686.6,0.0000,7592.2,4449.7,4252.8,3658.0,0.0000,-374.61,-115.05,-104.26,-44.932,-142.53,-587.69,0.0000,-1069.1,-1552.1,-750.73,-1231.7
1050.000000000,91.481,2035.1,2084.1,1929.3,312.81,4163.5,969.92,28.324,6359.3,2702.3,3360.2,2023.2,0.0000,-6675.5,-6930.6,-1430.8,-2230.3,-2253.7,-16007.,-117.26,-19611.,-6249.1,-4171.9,-2548.1,67.237,2395.3,2184.1,2032.9,343.44,4596.5,1686.6,0.0000,7592.2,4449.7,4252.8,3658.0,0.0000,-373.73,-114.78,-104.15,-44.825,-142.60,-587.69,0.0000,-1069.1,-1552.0,-750.72,-1231.6
1051.000000000,91.333,2031.3,2081.5,1929.2,312.17,4172.4,969.91,23.545,6360.4,2702.4,3360.2,2023.5,0.0000,-6676.2,-6930.8,-1432.1,-2229.7,-2256.7,-16005.,-117.21,-19611.,-6248.7,-4171.4,-2547.3,67.112,2390.8,2180.0,2032.4,342.85,4596.5,1686.6,0.0000,7592.2,4449.7,4252.8,3658.0,0.0000,-373.05,-114.57,-104.07,-44.741,-142.66,-587.69,0.0000,-1069.1,-1551.9,-750.71,-1231.5
1052.000000000,91.352,2027.3,2079.7,1928.6,311.69,4180.3,969.91,20.673,6370.2,2703.0,3360.1,2023.7,0.0000,-6676.6,-6930.9,-1433.3,-2229.1,-2259.9,-16004.,-117.15,-19611.,-6248.3,-4170.8,-2546.5,66.950,2385.1,2174.8,2031.6,342.09,4596.4,1686.6,0.0000,7592.2,4449.7,4252.8,3658.0,0.0000,-372.16,-114.30,-103.96,-44.633,-142.72,-587.69,0.0000,-1069.1,-1551.8,-750.69,-1231.3
1053.000000000,91.252,2024.3,2079.6,1928.1,311.06,4188.0,969.92,13.149,6370.5,2703.4,3360.1,2024.3,0.0000,-6677.0,-6930.8,-1434.4,-2228.5,-2263.7,-16003.,-117.10,-19610.,-6247.9,-4170.2,-2545.7,66.788,2379.3,2169.5,2030.9,341.34,4596.3,1686.6,0.0000,7592.2,4449.7,4252.8,3658.0,0.0000,-371.28,-114.03,-103.85,-44.526,-142.78,-587.69,0.0000,-1069.1,-1551.7,-750.68,-1231.2
1054.000000000,91.093,2020.1,2075.0,1927.4,310.44,4189.5,969.92,13.024,6370.3,2703.4,3360.1,2024.0,0.0000,-6677.2,-6930.5,-1435.4,-2227.9,-2267.1,-16001.,-117.04,-19610.,-6247.4,-4169.6,-2544.9,66.621,2373.3,2164.1,2030.1,340.56,4596.3,1686.6,0.0000,7592.2,4449.7,4252.8,3658.0,0.0000,-370.35,-113.74,-103.74,-44.414,-142.84,-587.69,0.0000,-1069.1,-1551.6,-750.66,-1231.1
1055.000000000,90.929,2015.4,2070.2,1927.2,309.82,4197.1,969.92,13.023,6370.0,2703.9,3360.0,2024.2,0.0000,-6677.1,-6930.0,-1436.3,-2227.3,-2270.2,-16000.,-116.98,-19610.,-6247.0,-4169.0,-2544.1,66.459,2367.6,2158.8,2029.4,339.80,4596.2,1686.6,0.0000,7592.2,4449.7,4252.8,3658.0,0.0000,-369.45,-113.46,-103.63,-44.306,-142.90,-587.69,0.0000,-1069.1,-1551.5,-750.65,-1231.0
1056.000000000,90.762,2010.8,2068.0,1927.9,309.18,4200.7,969.92,11.973,6369.7,2704.2,3360.0,2024.4,0.0000,-6676.8,-6929.5,-1437.2,-2226.6,-2273.0,-15998.,-116.93,-19609.,-6246.6,-4168.5,-2543.3,66.326,2362.8,2154.5,2028.8,339.18,4596.1,1686.6,0.0000,7592.2,4449.7,4252.8,3658.0,0.0000,-368.71,-113.23,-103.54,-44.217,-142.96,-587.69,0.0000,-1069.1,-1551.4,-750.64,-1230.9
1057.000000000,90.611,2006.6,2067.1,1927.2,308.60,4206.5,969.92,5.3942,6369.3,2704.4,3360.0,2024.6,0.0000,-6676.5,-6928.8,-1438.1,-2226.0,-2275.6,-15997.,-116.87,-19609.,-6246.2,-4167.9,-2542.5,66.193,2358.1,2150.2,2028.2,338.56,4596.1,1686.6,0.0000,7592.2,4449.7,4252.8,3658.0,0.0000,-367.97,-112.99,-103.45,-44.128,-143.01,-587.69,0.0000,-1069.1,-1551.3,-750.62,-1230.7
1058.000000000,90.463,2002.6,2063.9,1926.6,308.02,4209.6,969.92,5.4035,6368.9,2704.3,3360.0,2024.7,0.0000,-6676.0,-6928.1,-1438.9,-2225.3,-2278.0,-15995.,-116.82,-19609.,-6245.8,-4167.3,-2541.7,66.050,2353.0,2145.5,2027.6,337.89,4596.0,1686.6,0.0000,7592.2,4449.7,4252.8,3658.0,0.0000,-367.17,-112.74,-103.36,-44.033,-143.07,-587.69,0.0000,-1069.1,-1551.2,-750.61,-1230.6
1059.000000000,90.316,1998.4,2059.6,1926.0,307.45,4216.0,969.93,5.4042,6374.6,2704.0,3360.0,2024.7,0.0000,-6675.3,-6927.3,-1439.6,-2224.6,-2280.2,-15994.,-116.76,-19609.,-6245.4,-4166.7,-2540.9,65.887,2347.2,2140.2,2026.8,337.13,4596.0,1686.6,0.0000,7592.2,4449.7,4252.8,3658.0,0.0000,-366.25,-112.45,-103.25,-43.925,-143.12,-587.69,0.0000,-1069.1,-1551.1,-750.59,-1230.5
1060.000000000,90.161,1994.0,2055.3,1925.5,306.85,4215.4,969.92,5.4048,6379.1,2704.0,3359.9,2024.7,0.0000,-6674.4,-6926.3,-1440.4,-2223.9,-2282.4,-15992.,-116.70,-19610.,-6244.9,-4166.1,-2540.1,65.750,2342.3,2135.8,2026.2,336.50,4595.9,1686.6,0.0000,7592.2,4449.7,4252.8,3658.0,0.0000,-365.48,-112.21,-103.16,-43.834,-143.17,-587.69,0.0000,-1069.1,-1551.0,-750.58,-1230.4
1061.000000000,90.017,1990.2,2052.4,1925.0,306.39,4220.4,969.88,5.4054,6380.9,2704.0,3360.0,2024.8,0.0000,-6673.4,-6925.4,-1441.0,-2223.2,-2284.4,-15991.,-116.65,-19610.,-6244.5,-4165.6,-2539.3,65.735,2341.8,2135.3,2026.2,341.21,4595.9,1686.6,0.0000,7592.2,4449.7,4264.6,3684.5,0.0000,-365.38,-112.17,-103.15,-43.853,-143.22,-587.69,0.0000,-1069.1,-1550.9,-750.62,-1230.9
1062.000000000,89.944,1994.0,2055.8,1924.3,307.16,4224.7,969.88,5.4059,6383.8,2703.9,3360.1,2024.8,0.0000,-6672.8,-6924.7,-1441.7,-2222.5,-2286.4,-15989.,-116.59,-19610.,-6244.1,-4165.0,-2538.5,459.76,2751.4,2663.2,2083.4,403.22,4634.7,1686.6,438.98,7692.1,4586.9,4373.3,3818.9,0.0000,-372.97,-124.71,-103.99,-45.039,-143.45,-587.69,-20.055,-1070.6,-1550.8,-751.17,-1234.1
1063.000000000,90.555,2010.1,2069.2,1924.1,309.70,4224.3,969.89,5.4066,6383.6,2703.8,3360.2,2024.9,0.0000,-6673.4,-6924.8,-1442.4,-2222.0,-2288.2,-15988.,-116.54,-19610.,-6243.7,-4164.4,-2537.8,67.485,2404.1,2192.1,2034.3,344.59,4596.7,1686.6,0.0000,7592.6,4450.0,4252.9,3658.0,0.0000,-375.10,-115.16,-104.31,-44.990,-143.32,-587.69,0.0000,-1069.2,-1550.7,-750.53,-1230.0
1064.000000000,90.911,2022.4,2081.8,1925.4,311.11,4224.1,969.89,5.4072,6384.6,2703.7,3360.2,2025.0,0.0000,-6674.7,-6925.3,-1443.1,-2221.6,-2290.0,-15987.,-116.49,-19609.,-6243.2,-4163.9,-2537.0,67.579,2407.5,2195.2,2034.5,345.03,4596.6,1686.6,0.0000,7592.2,4449.7,4252.8,3658.0,0.0000,-375.63,-115.32,-104.38,-45.052,-143.36,-587.69,0.0000,-1069.2,-1550.6,-750.52,-1229.9
1065.000000000,91.114,2028.1,2087.7,1926.6,312.64,4224.0,969.89,5.4078,6394.0,2703.7,3360.2,2025.1,0.0000,-6676.1,-6925.9,-1443.8,-2221.1,-2291.7,-15985.,-116.43,-19609.,-6242.8,-4163.3,-2536.2,67.571,2407.2,2195.0,2034.4,344.99,4596.6,1686.6,0.0000,7592.2,4449.7,4252.8,3658.0,0.0000,-375.59,-115.32,-104.37,-45.047,-143.41,-587.69,0.0000,-1069.2,-1550.5,-750.50,-1229.7
1066.000000000,91.406,2030.2,2090.1,1926.9,313.20,4223.7,969.86,5.4084,6397.9,2703.7,3360.2,2025.2,0.0000,-6677.4,-6926.3,-1444.4,-2220.7,-2293.3,-15984.,-116.38,-19609.,-6242.4,-4162.7,-2535.4,67.519,2405.3,2193.3,2034.2,344.75,4596.5,1686.6,0.0000,7592.2,4449.7,4252.8,3658.0,0.0000,-375.31,-115.24,-104.34,-45.013,-143.45,-587.69,0.0000,-1069.2,-1550.4,-750.49,-1229.6
1067.000000000,91.460,2030.3,2090.6,1926.7,313.16,4223.3,969.85,5.4090,6399.0,2703.6,3360.2,2025.4,0.0000,-6678.4,-6926.5,-1445.0,-2220.1,-2294.9,-15982.,-116.32,-19608.,-6241.9,-4162.2,-2534.6,67.441,2402.5,2190.7,2033.8,344.38,4596.5,1686.6,0.0000,7592.1,4449.7,4252.8,3658.0,0.0000,-374.88,-115.11,-104.28,-44.960,-143.50,-587.69,0.0000,-1069.2,-1550.3,-750.48,-1229.5
1068.000000000,91.342,2029.3,2089.8,1926.7,312.92,4223.0,969.85,5.4095,6398.9,2704.0,3360.2,2025.5,0.0000,-6679.0,-6926.6,-1445.6,-2219.6,-2296.4,-15981.,-116.27,-19608.,-6241.5,-4161.6,-2533.8,67.344,2399.1,2187.6,2033.4,343.93,4596.5,1686.6,0.0000,7592.1,4449.7,4252.8,3658.0,0.0000,-374.35,-114.95,-104.22,-44.896,-143.54,-587.69,0.0000,-1069.2,-1550.2,-750.46,-1229.4
1069.000000000,91.272,2027.3,2088.6,1929.9,312.57,4222.6,969.85,5.4101,6398.7,2704.1,3360.2,2025.6,0.0000,-6679.5,-6926.5,-1446.1,-2219.0,-2297.8,-15979.,-116.21,-19607.,-6241.0,-4161.1,-2533.0,67.235,2395.2,2184.0,2032.9,343.43,4596.4,1686.6,0.0000,7592.1,4449.7,4252.8,3658.0,0.0000,-373.75,-114.76,-104.15,-44.824,-143.58,-587.69,0.0000,-1069.2,-1550.1,-750.45,-1229.3
1070.000000000,91.203,2025.9,2087.3,1931.1,312.17,4222.2,969.85,5.4161,6398.6,2704.1,3360.2,2025.6,0.0000,-6679.8,-6926.3,-1446.6,-2218.4,-2299.2,-15978.,-116.16,-19607.,-6240.6,-4160.5,-2532.2,67.118,2391.1,2180.2,2032.3,342.88,4596.4,1686.6,0.0000,7592.1,4449.7,4252.8,3658.0,0.0000,-373.10,-114.56,-104.07,-44.746,-143.62,-587.69,0.0000,-1069.2,-1550.0,-750.43,-1229.1
1071.000000000,91.092,2023.4,2084.9,1931.2,311.74,4221.8,969.85,5.4236,6398.5,2704.1,3360.2,2025.7,0.0000,-6679.8,-6926.0,-1447.0,-2217.8,-2300.5,-15976.,-116.10,-19606.,-6240.1,-4159.9,-2531.4,66.996,2386.7,2176.3,2031.8,342.31,4596.4,1686.6,0.0000,7592.1,4449.7,4252.8,3658.0,0.0000,-372.42,-114.35,-103.99,-44.664,-143.66,-587.69,0.0000,-1069.2,-1549.9,-750.42,-1229.0
1072.000000000,90.972,2020.3,2081.9,1931.1,311.25,4221.0,969.85,5.4288,6398.3,2704.4,3360.2,2025.8,0.0000,-6679.6,-6925.6,-1447.4,-2217.2,-2301.7,-15975.,-116.05,-19605.,-6239.7,-4159.4,-2530.6,66.866,2382.1,2172.0,2028.4,341.65,4589.0,1686.6,0.0000,7587.7,4449.7,4252.8,3658.0,0.0000,-371.69,-114.13,-103.80,-44.577,-143.47,-587.69,0.0000,-1069.1,-1549.8,-750.40,-1228.9
1073.000000000,90.844,2017.7,2078.7,1932.0,310.72,4218.0,969.86,5.4369,6397.7,2704.9,3360.2,2026.0,0.0000,-6679.1,-6925.1,-1447.7,-2216.5,-2302.8,-15974.,-115.99,-19604.,-6239.2,-4158.8,-2529.8,66.725,2377.0,2167.5,2018.4,340.84,4564.6,1686.6,0.0000,7572.9,4449.7,4252.8,3658.0,0.0000,-370.90,-113.88,-103.39,-44.483,-142.72,-587.69,0.0000,-1069.0,-1549.7,-750.39,-1228.8
1074.000000000,90.708,2014.5,2075.4,1930.7,310.05,4210.8,969.86,5.4327,6396.0,2705.3,3360.1,2026.2,0.0000,-6678.3,-6924.5,-1447.9,-2215.8,-2303.7,-15972.,-115.94,-19604.,-6238.8,-4158.3,-2529.0,66.579,2371.9,2162.7,2008.3,339.99,4540.0,1686.6,0.0000,7558.0,4449.7,4252.8,3658.0,0.0000,-370.08,-113.63,-102.97,-44.386,-141.97,-587.69,0.0000,-1068.9,-1549.6,-750.37,-1228.6
1075.000000000,90.564,2010.6,2071.6,1924.7,309.30,4200.3,969.86,5.4269,6392.9,2705.3,3360.2,2026.3,0.0000,-6677.3,-6923.9,-1447.8,-2215.2,-2304.3,-15971.,-115.88,-19603.,-6238.4,-4157.7,-2528.3,66.429,2366.5,2157.9,1998.1,339.13,4515.2,1686.6,0.0000,7542.9,4449.7,4252.8,3658.0,0.0000,-369.24,-113.36,-102.54,-44.286,-141.20,-587.69,0.0000,-1068.8,-1549.5,-750.36,-1228.5
1076.000000000,90.415,2008.3,2067.9,1917.1,308.55,4190.3,969.86,5.4274,6388.8,2705.3,3360.3,2026.4,0.0000,-6676.1,-6923.1,-1447.6,-2214.5,-2304.6,-15969.,-115.83,-19602.,-6237.9,-4157.2,-2527.5,66.278,2361.1,2152.9,1987.9,338.26,4490.5,1686.6,0.0000,7527.9,4449.7,4252.8,3658.0,0.0000,-368.38,-113.09,-102.12,-44.185,-140.43,-587.69,0.0000,-1068.7,-1549.4,-750.35,-1228.4
1077.000000000,90.275,2010.9,2070.5,1910.0,308.92,4182.9,969.86,5.4280,6384.0,2705.0,3360.3,2026.4,0.0000,-6675.4,-6922.6,-1447.4,-2213.8,-2304.8,-15968.,-115.77,-19601.,-6237.5,-4156.6,-2526.7,371.79,2736.3,2675.4,2057.0,391.90,4571.7,1686.6,347.11,7632.9,4542.6,4335.8,3774.4,0.0000,-375.87,-125.50,-103.56,-45.312,-142.09,-587.69,-15.856,-1070.0,-1549.3,-750.76,-1231.1
1078.000000000,90.864,2026.5,2082.8,1908.3,311.41,4180.7,969.86,5.4286,6379.6,2705.4,3360.3,2026.5,0.0000,-6675.8,-6922.8,-1447.3,-2213.3,-2305.1,-15966.,-115.72,-19600.,-6237.1,-4156.1,-2525.9,67.946,2420.5,2207.1,2006.7,346.87,4521.0,1686.6,0.0000,7546.3,4450.8,4256.2,3659.8,0.0000,-377.65,-115.94,-103.59,-45.301,-141.36,-587.69,0.0000,-1068.9,-1549.3,-750.34,-1228.2
1079.000000000,91.201,2038.1,2094.1,1908.1,312.61,4175.4,969.86,5.4292,6374.0,2705.5,3360.5,2026.6,0.0000,-6676.9,-6923.4,-1447.2,-2212.8,-2305.7,-15965.,-115.67,-19599.,-6236.7,-4155.5,-2525.1,68.007,2422.7,2209.1,1997.5,346.59,4497.0,1686.6,0.0000,7531.1,4449.9,4255.0,3658.9,0.0000,-377.99,-116.05,-103.33,-45.339,-140.64,-587.69,0.0000,-1068.7,-1549.2,-750.31,-1228.1
1080.000000000,91.496,2043.0,2098.9,1906.9,313.88,4163.5,969.86,5.4297,6366.0,2705.3,3360.5,2026.7,0.0000,-6678.0,-6924.0,-1447.0,-2212.4,-2306.0,-15963.,-115.61,-19598.,-6236.2,-4155.0,-2524.3,67.988,2422.0,2208.5,1988.5,346.25,4473.5,1686.6,0.0000,7516.9,4449.8,4254.1,3658.5,0.0000,-377.90,-116.03,-103.01,-45.326,-139.91,-587.69,0.0000,-1068.6,-1549.1,-750.30,-1227.9
1081.000000000,91.610,2044.3,2101.0,1902.1,314.13,4149.0,969.86,5.4344,6358.0,2705.5,3360.6,2026.8,0.0000,-6679.0,-6924.4,-1446.9,-2211.9,-2306.0,-15962.,-115.56,-19597.,-6235.8,-4154.4,-2523.5,67.937,2420.2,2206.8,1979.5,345.78,4450.4,1686.6,0.0000,7502.9,4449.7,4253.4,3658.2,0.0000,-377.62,-115.95,-102.68,-45.292,-139.20,-587.69,0.0000,-1068.5,-1549.0,-750.28,-1227.8
1082.000000000,91.511,2044.1,2101.2,1895.6,313.90,4133.0,969.86,5.4482,6355.9,2706.3,3360.5,2026.9,0.0000,-6679.8,-6924.6,-1446.5,-2211.4,-2305.8,-15960.,-115.50,-19596.,-6235.3,-4153.9,-2522.8,67.861,2417.5,2204.4,1970.5,345.25,4427.6,1686.6,0.0000,7489.2,4449.7,4253.1,3658.0,0.0000,-377.21,-115.82,-102.33,-45.241,-138.48,-587.69,0.0000,-1068.4,-1548.9,-750.26,-1227.7
1083.000000000,91.463,2042.9,2100.2,1887.9,313.50,4121.4,969.86,5.4522,6353.6,2706.7,3360.3,2027.1,0.0000,-6680.3,-6924.8,-1445.9,-2210.8,-2305.4,-15959.,-115.45,-19595.,-6234.9,-4153.4,-2522.0,67.768,2414.2,2201.4,1961.4,344.65,4404.8,1686.6,0.0000,7475.4,4449.7,4252.9,3658.0,0.0000,-376.70,-115.67,-101.97,-45.179,-137.76,-587.69,0.0000,-1068.3,-1548.8,-750.25,-1227.6
1084.000000000,91.386,2040.7,2099.4,1884.1,313.01,4109.6,969.73,5.4527,6347.1,2706.5,3360.2,2027.2,0.0000,-6680.5,-6924.7,-1445.2,-2210.2,-2304.8,-15957.,-115.40,-19594.,-6234.5,-4152.8,-2521.2,67.654,2410.1,2197.6,1951.9,343.96,4381.5,1686.6,0.0000,7461.3,4449.7,4252.8,3658.0,0.0000,-376.06,-115.48,-101.59,-45.103,-137.01,-587.69,0.0000,-1068.2,-1548.7,-750.23,-1227.4
1085.000000000,91.286,2039.0,2098.4,1877.2,312.43,4092.3,969.69,5.4533,6337.9,2706.2,3360.2,2027.3,0.0000,-6680.7,-6924.6,-1444.4,-2209.6,-2304.1,-15956.,-115.34,-19593.,-6234.1,-4152.3,-2520.4,67.521,2405.4,2193.3,1942.2,343.19,4357.8,1686.6,0.0000,7446.9,4449.7,4252.8,3658.0,0.0000,-375.32,-115.25,-101.19,-45.014,-136.25,-587.69,0.0000,-1068.1,-1548.6,-750.22,-1227.3
1086.000000000,91.167,2036.3,2096.4,1869.4,311.78,4072.8,969.69,5.4538,6327.2,2706.2,3360.3,2027.4,0.0000,-6680.6,-6924.3,-1443.5,-2209.0,-2303.2,-15954.,-115.29,-19591.,-6233.6,-4151.7,-2519.6,67.384,2400.5,2188.9,1932.6,342.39,4334.2,1686.6,0.0000,7432.6,4449.7,4252.8,3658.0,0.0000,-374.56,-115.01,-100.79,-44.923,-135.49,-587.69,0.0000,-1068.0,-1548.5,-750.21,-1227.2
1087.000000000,91.037,2033.1,2092.8,1861.1,311.08,4053.1,969.67,5.4544,6315.6,2706.2,3360.5,2027.5,0.0000,-6680.2,-6923.8,-1442.5,-2208.3,-2302.1,-15953.,-115.23,-19590.,-6233.2,-4151.2,-2518.8,67.239,2395.3,2184.2,1922.8,341.56,4310.4,1686.6,0.0000,7418.2,4449.7,4252.8,3658.0,0.0000,-373.75,-114.76,-100.38,-44.826,-134.71,-587.69,0.0000,-1067.9,-1548.4,-750.19,-1227.1
1088.000000000,90.895,2030.1,2089.2,1852.5,310.35,4034.3,969.66,5.4601,6304.5,2706.2,3360.6,2027.7,0.0000,-6679.6,-6923.2,-1441.4,-2207.7,-2301.0,-15951.,-115.18,-19589.,-6232.7,-4150.7,-2518.0,67.087,2389.9,2179.2,1913.0,340.69,4286.5,1686.6,0.0000,7403.7,4449.7,4252.8,3658.0,0.0000,-372.90,-114.49,-99.964,-44.725,-133.93,-587.69,0.0000,-1067.8,-1548.3,-750.18,-1226.9
1089.000000000,90.745,2026.4,2086.2,1843.9,309.60,4017.8,969.66,5.4690,6293.3,2706.3,3360.6,2027.8,0.0000,-6678.7,-6922.6,-1440.2,-2207.0,-2299.6,-15950.,-115.12,-19588.,-6232.3,-4150.1,-2517.3,66.934,2384.5,2174.2,1903.1,339.82,4262.8,1686.6,0.0000,7389.3,4449.7,4252.8,3658.0,0.0000,-372.04,-114.22,-99.549,-44.622,-133.15,-587.69,0.0000,-1067.6,-1548.2,-750.17,-1226.8
1090.000000000,90.592,2022.2,2082.8,1835.3,308.84,4000.6,969.67,5.4696,6281.2,2706.3,3360.6,2027.9,0.0000,-6677.6,-6921.8,-1438.9,-2206.3,-2298.2,-15948.,-115.07,-19586.,-6231.8,-4149.6,-2516.5,66.784,2379.1,2169.4,1893.5,338.97,4239.4,1686.6,0.0000,7375.1,4449.7,4252.8,3658.0,0.0000,-371.19,-113.96,-99.141,-44.523,-132.38,-587.69,0.0000,-1067.5,-1548.1,-750.15,-1226.7
1091.000000000,90.450,2024.3,2084.6,1827.2,309.09,3982.7,969.67,5.4701,6269.7,2706.4,3360.5,2028.0,0.0000,-6676.8,-6921.3,-1437.8,-2205.7,-2296.7,-15947.,-115.02,-19585.,-6231.4,-4149.0,-2515.7,322.32,2653.5,2576.7,1954.4,391.93,4312.8,1686.6,267.81,7464.7,4529.8,4338.0,3760.8,0.0000,-377.62,-123.75,-100.26,-45.543,-133.51,-587.69,-12.232,-1068.7,-1548.0,-750.58,-1229.0
1092.000000000,90.954,2037.3,2095.6,1823.5,311.16,3971.9,969.67,5.4826,6259.9,2706.3,3360.5,2028.1,0.0000,-6677.1,-6921.4,-1436.7,-2205.1,-2295.3,-15945.,-114.96,-19583.,-6231.0,-4148.5,-2514.9,129.78,2495.9,2295.8,1937.5,380.35,4287.9,1686.6,64.246,7428.2,4495.3,4295.2,3702.8,0.0000,-379.40,-118.14,-100.40,-45.708,-133.14,-587.69,-2.9345,-1068.2,-1548.0,-750.34,-1227.5
1093.000000000,91.355,2048.6,2106.8,1822.3,312.42,3965.8,969.67,5.4882,6251.2,2706.3,3360.5,2028.2,0.0000,-6678.1,-6921.9,-1435.8,-2204.7,-2294.2,-15944.,-114.91,-19582.,-6230.5,-4148.0,-2514.2,68.543,2441.8,2226.5,1902.6,347.25,4243.5,1686.6,0.0000,7377.2,4449.7,4253.0,3658.0,0.0000,-380.97,-116.97,-100.36,-45.695,-132.41,-587.69,0.0000,-1067.5,-1547.9,-750.11,-1226.3
1094.000000000,91.823,2056.6,2114.2,1820.7,314.10,3955.4,969.67,5.5020,6241.7,2706.5,3360.7,2028.4,0.0000,-6679.4,-6922.5,-1434.9,-2204.2,-2292.9,-15942.,-114.86,-19581.,-6230.1,-4147.4,-2513.4,68.606,2444.0,2228.6,1895.1,347.41,4223.1,1686.6,0.0000,7364.8,4449.7,4253.0,3658.0,0.0000,-381.33,-117.08,-100.13,-45.738,-131.73,-587.69,0.0000,-1067.4,-1547.8,-750.10,-1226.2
1095.000000000,92.178,2060.2,2118.4,1816.8,314.60,3941.2,969.67,5.5025,6232.5,2706.6,3360.6,2028.5,0.0000,-6680.6,-6923.1,-1434.0,-2203.8,-2291.5,-15941.,-114.81,-19579.,-6229.6,-4146.9,-2512.6,68.584,2443.3,2227.9,1886.9,347.17,4202.1,1686.6,0.0000,7352.0,4449.7,4252.9,3658.0,0.0000,-381.22,-117.06,-99.840,-45.723,-131.03,-587.69,0.0000,-1067.3,-1547.7,-750.08,-1226.1
1096.000000000,92.308,2061.1,2119.6,1811.7,314.69,3924.4,969.66,5.5031,6224.7,2706.8,3360.6,2028.6,0.0000,-6681.7,-6923.5,-1433.0,-2203.3,-2289.8,-15939.,-114.75,-19577.,-6229.2,-4146.4,-2511.8,68.521,2441.0,2225.8,1878.5,346.70,4180.8,1686.6,0.0000,7339.1,4449.7,4252.8,3658.0,0.0000,-380.87,-116.95,-99.519,-45.681,-130.33,-587.69,0.0000,-1067.2,-1547.6,-750.07,-1226.0
1097.000000000,92.325,2060.9,2119.3,1805.0,314.44,3910.4,969.63,5.5036,6219.4,2707.1,3360.7,2028.7,0.0000,-6682.5,-6923.8,-1431.9,-2202.7,-2288.0,-15937.,-114.70,-19576.,-6228.7,-4145.8,-2511.1,68.441,2438.2,2223.2,1870.2,346.18,4160.2,1686.6,0.0000,7326.6,4449.7,4252.8,3658.0,0.0000,-380.44,-116.82,-99.194,-45.627,-129.63,-587.69,0.0000,-1067.1,-1547.5,-750.06,-1225.9
1098.000000000,92.630,2060.5,2119.6,1797.6,314.20,3898.4,969.64,5.5051,6213.6,2707.2,3360.8,2028.9,0.0000,-6683.1,-6924.0,-1430.7,-2202.2,-2286.1,-15936.,-114.65,-19574.,-6228.3,-4145.3,-2510.3,68.548,2442.0,2226.7,1865.5,346.59,4146.8,1686.6,0.0000,7318.5,4449.7,4252.8,3658.0,0.0000,-381.04,-117.01,-99.089,-45.699,-129.17,-587.69,0.0000,-1067.0,-1547.4,-750.04,-1225.7
1099.000000000,92.969,2061.6,2121.0,1791.1,314.09,3884.6,969.64,5.5205,6205.5,2707.2,3360.8,2029.0,0.0000,-6683.8,-6924.1,-1429.4,-2201.6,-2284.1,-15934.,-114.59,-19573.,-6227.8,-4144.7,-2509.5,68.437,2438.0,2223.1,1857.0,345.93,4126.0,1686.6,0.0000,7305.8,4449.7,4252.8,3658.0,0.0000,-380.43,-116.83,-98.741,-45.625,-128.47,-587.69,0.0000,-1066.9,-1547.3,-750.03,-1225.6
1100.000000000,92.932,2060.6,2121.2,1785.3,313.64,3868.5,969.64,5.5211,6195.7,2707.2,3360.8,2029.2,0.0000,-6684.2,-6924.1,-1428.1,-2201.1,-2282.1,-15933.,-114.54,-19571.,-6227.4,-4144.2,-2508.7,68.317,2433.8,2219.2,1848.5,345.23,4105.1,1686.6,0.0000,7293.2,4449.7,4252.8,3658.0,0.0000,-379.77,-116.62,-98.387,-45.545,-127.76,-587.69,0.0000,-1066.8,-1547.2,-750.01,-1225.5
1101.000000000,92.860,2058.6,2119.3,1778.8,313.22,3850.4,969.64,5.5230,6184.7,2707.6,3360.8,2029.3,0.0000,-6684.4,-6923.9,-1426.7,-2200.5,-2279.9,-15931.,-114.49,-19570.,-6227.0,-4143.7,-2507.9,68.184,2429.0,2214.8,1839.8,344.47,4084.0,1686.6,0.0000,7280.4,4449.7,4252.8,3658.0,0.0000,-379.03,-116.40,-98.020,-45.456,-127.04,-587.69,0.0000,-1066.7,-1547.1,-750.00,-1225.4
1102.000000000,92.759,2056.5,2116.5,1771.3,312.56,3832.5,969.64,5.5314,6173.4,2707.4,3360.7,2029.5,0.0000,-6684.3,-6923.6,-1425.3,-2199.9,-2277.6,-15929.,-114.43,-19568.,-6226.6,-4143.1,-2507.2,68.039,2423.9,2210.2,1830.9,343.66,4062.6,1686.6,0.0000,7267.4,4449.7,4252.8,3658.0,0.0000,-378.23,-116.15,-97.643,-45.360,-126.32,-587.69,0.0000,-1066.6,-1547.0,-749.99,-1225.2
1103.000000000,92.667,2053.3,2113.4,1763.7,311.86,3814.6,969.62,5.5268,6162.9,2707.3,3360.8,2029.7,0.0000,-6684.0,-6923.2,-1423.8,-2199.2,-2275.2,-15928.,-114.38,-19566.,-6226.1,-4142.6,-2506.4,67.886,2418.4,2205.2,1821.9,342.80,4041.0,1686.6,0.0000,7254.3,4449.7,4252.8,3658.0,0.0000,-377.38,-115.88,-97.256,-45.258,-125.58,-587.69,0.0000,-1066.4,-1547.0,-749.97,-1225.1
1104.000000000,92.522,2049.7,2110.3,1756.2,311.05,3797.1,969.60,5.5271,6152.5,2707.5,3360.8,2029.7,0.0000,-6683.3,-6922.7,-1422.2,-2198.6,-2272.7,-15926.,-114.33,-19564.,-6225.7,-4142.1,-2505.6,67.735,2413.0,2200.3,1813.0,341.95,4019.6,1686.6,0.0000,7241.3,4449.7,4252.8,3658.0,0.0000,-376.53,-115.62,-96.874,-45.157,-124.85,-587.69,0.0000,-1066.3,-1546.9,-749.96,-1225.0
1105.000000000,92.371,2045.8,2107.4,1748.2,310.32,3779.1,969.58,5.5276,6141.5,2707.6,3360.9,2029.9,0.0000,-6682.5,-6922.1,-1420.6,-2197.9,-2270.1,-15925.,-114.27,-19563.,-6225.2,-4141.5,-2504.9,67.611,2408.6,2196.2,1804.8,341.24,3999.7,1686.6,0.0000,7229.2,4449.7,4252.8,3658.0,0.0000,-375.83,-115.40,-96.529,-45.074,-124.16,-587.69,0.0000,-1066.2,-1546.8,-749.95,-1224.9
1106.000000000,92.230,2042.4,2104.5,1740.2,309.65,3760.9,969.58,5.5281,6130.6,2707.7,3361.2,2030.0,0.0000,-6681.6,-6921.4,-1418.9,-2197.2,-2267.5,-15923.,-114.22,-19561.,-6224.8,-4141.0,-2504.1,67.484,2404.1,2192.1,1796.6,340.52,3979.8,1686.6,0.0000,7217.2,4449.7,4252.8,3658.0,0.0000,-375.11,-115.17,-96.184,-44.990,-123.47,-587.69,0.0000,-1066.1,-1546.7,-749.93,-1224.7
1107.000000000,92.092,2039.1,2101.0,1732.5,308.98,3742.5,969.58,5.5287,6119.3,2707.8,3361.4,2030.2,0.0000,-6680.5,-6920.7,-1417.2,-2196.6,-2264.8,-15921.,-114.17,-19559.,-6224.4,-4140.5,-2503.3,67.353,2399.4,2187.9,1788.4,339.78,3959.9,1686.6,0.0000,7205.0,4449.7,4252.8,3658.0,0.0000,-374.37,-114.94,-95.834,-44.902,-122.78,-587.69,0.0000,-1066.0,-1546.6,-749.92,-1224.6
1108.000000000,91.956,2035.8,2097.1,1724.7,308.32,3724.0,969.58,5.5292,6107.8,2708.0,3361.3,2030.3,0.0000,-6679.3,-6919.9,-1415.5,-2195.9,-2262.0,-15920.,-114.11,-19557.,-6223.9,-4139.9,-2502.5,67.213,2394.4,2183.3,1780.0,338.99,3939.6,1686.6,0.0000,7192.8,4449.7,4252.8,3658.0,0.0000,-373.58,-114.69,-95.474,-44.809,-122.08,-587.69,0.0000,-1065.9,-1546.5,-749.91,-1224.5
1109.000000000,91.961,2032.2,2093.1,1717.0,307.66,3705.7,969.58,5.5297,6096.7,2708.0,3361.3,2030.4,0.0000,-6677.8,-6919.0,-1413.7,-2195.1,-2259.2,-15918.,-114.06,-19556.,-6223.5,-4139.4,-2501.8,67.066,2389.2,2178.6,1771.5,338.17,3919.1,1686.6,0.0000,7180.3,4449.7,4252.8,3658.0,0.0000,-372.74,-114.42,-95.107,-44.711,-121.37,-587.69,0.0000,-1065.8,-1546.4,-749.89,-1224.4
1110.000000000,91.957,2028.1,2089.1,1709.3,306.98,3687.4,969.58,5.5303,6085.7,2708.0,3361.1,2030.5,0.0000,-6676.2,-6918.1,-1411.9,-2194.4,-2256.3,-15916.,-114.01,-19554.,-6223.1,-4138.9,-2501.0,66.911,2383.7,2173.5,1762.8,337.32,3898.4,1686.6,0.0000,7167.8,4449.7,4252.8,3658.0,0.0000,-371.86,-114.14,-94.731,-44.608,-120.64,-587.69,0.0000,-1065.6,-1546.3,-749.88,-1224.3
1111.000000000,91.654,2023.8,2084.8,1701.4,306.24,3668.8,969.58,5.5308,6075.0,2708.1,3360.9,2030.6,0.0000,-6674.3,-6917.1,-1410.0,-2193.7,-2253.3,-15915.,-113.96,-19552.,-6222.6,-4138.3,-2500.2,66.755,2378.1,2168.4,1754.1,336.45,3877.6,1686.6,0.0000,7155.2,4449.7,4252.8,3658.0,0.0000,-370.97,-113.86,-94.354,-44.503,-119.92,-587.69,0.0000,-1065.5,-1546.2,-749.87,-1224.1
1112.000000000,91.317,2019.5,2080.7,1693.5,305.50,3653.2,969.58,5.5313,6063.8,2708.6,3360.8,2030.7,0.0000,-6672.3,-6915.9,-1408.2,-2192.9,-2250.3,-15913.,-113.90,-19550.,-6222.2,-4137.8,-2499.5,66.619,2373.3,2164.0,1746.0,335.69,3858.0,1686.6,0.0000,7143.2,4449.7,4252.8,3658.0,0.0000,-370.19,-113.61,-94.005,-44.413,-119.23,-587.69,0.0000,-1065.4,-1546.1,-749.85,-1224.0
1113.000000000,91.170,2015.4,2076.5,1685.9,304.79,3637.3,969.58,5.5318,6052.8,2708.9,3360.8,2030.8,0.0000,-6670.2,-6914.8,-1406.2,-2192.2,-2247.2,-15911.,-113.85,-19548.,-6221.8,-4137.3,-2498.7,66.484,2368.4,2159.6,1737.9,334.92,3838.4,1686.6,0.0000,7131.4,4449.7,4252.8,3658.0,0.0000,-369.41,-113.36,-93.657,-44.323,-118.54,-587.69,0.0000,-1065.3,-1546.1,-749.84,-1223.9
1114.000000000,91.023,2011.5,2072.5,1678.0,304.10,3619.3,969.58,5.5364,6041.6,2708.7,3360.8,2030.9,0.0000,-6667.9,-6913.5,-1404.3,-2191.4,-2244.0,-15909.,-113.80,-19546.,-6221.4,-4136.7,-2497.9,66.343,2363.4,2155.1,1729.7,334.14,3818.7,1686.6,0.0000,7119.4,4449.7,4252.8,3658.0,0.0000,-368.60,-113.10,-93.304,-44.229,-117.84,-587.69,0.0000,-1065.2,-1546.0,-749.83,-1223.8
1115.000000000,90.878,2007.3,2068.7,1670.2,303.42,3601.3,969.59,5.5452,6030.3,2708.6,3361.0,2031.1,0.0000,-6665.6,-6912.3,-1402.3,-2190.6,-2240.9,-15908.,-113.74,-19544.,-6221.0,-4136.2,-2497.1,66.190,2358.0,2150.1,1721.2,333.29,3798.5,1686.6,0.0000,7107.2,4449.7,4252.8,3658.0,0.0000,-367.71,-112.82,-92.936,-44.127,-117.13,-587.69,0.0000,-1065.1,-1545.9,-749.81,-1223.6
1116.000000000,90.640,2003.0,2064.4,1662.4,302.70,3583.1,969.59,5.5458,6018.9,2709.0,3360.9,2031.1,0.0000,-6663.1,-6910.9,-1400.3,-2189.8,-2237.6,-15906.,-113.69,-19542.,-6220.6,-4135.6,-2496.4,66.041,2352.7,2145.3,1712.9,332.47,3778.6,1686.6,0.0000,7095.1,4449.7,4252.8,3658.0,0.0000,-366.85,-112.54,-92.575,-44.027,-116.43,-587.69,0.0000,-1064.9,-1545.8,-749.80,-1223.5
1117.000000000,90.301,1998.7,2060.1,1654.8,301.98,3565.1,969.59,5.5463,6007.5,2709.2,3360.8,2031.2,0.0000,-6660.5,-6909.5,-1398.3,-2189.0,-2234.3,-15904.,-113.64,-19540.,-6220.2,-4135.1,-2495.6,65.899,2347.6,2140.6,1704.8,331.68,3759.1,1686.6,0.0000,7083.2,4449.7,4252.8,3658.0,0.0000,-366.03,-112.28,-92.224,-43.933,-115.74,-587.69,0.0000,-1064.8,-1545.7,-749.78,-1223.4
1118.000000000,90.234,1994.5,2056.4,1647.2,301.27,3547.1,969.59,5.5468,5996.4,2709.1,3360.7,2031.5,0.0000,-6657.9,-6908.1,-1396.3,-2188.2,-2230.9,-15903.,-113.59,-19538.,-6219.8,-4134.6,-2494.8,65.766,2342.9,2136.3,1696.9,330.93,3740.0,1686.6,0.0000,7071.7,4449.7,4252.8,3658.0,0.0000,-365.25,-112.03,-91.885,-43.844,-115.06,-587.69,0.0000,-1064.7,-1545.6,-749.77,-1223.3
1119.000000000,90.230,1990.4,2052.8,1639.6,300.59,3529.6,969.59,5.5473,5985.3,2708.5,3360.8,2031.7,0.0000,-6655.1,-6906.6,-1394.2,-2187.4,-2227.6,-15901.,-113.54,-19536.,-6219.3,-4134.0,-2494.0,65.631,2338.1,2131.9,1689.0,330.18,3721.1,1686.6,0.0000,7060.2,4449.7,4252.8,3658.0,0.0000,-364.47,-111.77,-91.546,-43.754,-114.38,-587.69,0.0000,-1064.6,-1545.5,-749.76,-1223.1
1120.000000000,90.124,1986.5,2048.9,1631.9,299.90,3511.9,969.59,5.5478,5974.4,2708.3,3360.8,2031.8,0.0000,-6652.3,-6905.1,-1392.1,-2186.6,-2224.1,-15899.,-113.48,-19534.,-6218.9,-4133.5,-2493.3,65.479,2332.7,2127.0,1680.8,329.34,3701.4,1686.6,0.0000,7048.2,4449.7,4252.8,3658.0,0.0000,-363.58,-111.49,-91.186,-43.653,-113.68,-587.69,0.0000,-1064.5,-1545.4,-749.74,-1223.0
1121.000000000,89.975,1982.4,2044.7,1624.2,299.19,3494.4,969.59,5.5483,5963.4,2708.2,3360.8,2031.9,0.0000,-6649.3,-6903.6,-1390.0,-2185.8,-2220.7,-15897.,-113.43,-19532.,-6218.5,-4132.9,-2492.5,65.324,2327.1,2122.0,1672.5,328.48,3681.6,1686.6,0.0000,7036.2,4449.7,4252.8,3658.0,0.0000,-362.68,-111.20,-90.822,-43.549,-112.97,-587.69,0.0000,-1064.4,-1545.3,-749.73,-1222.9
1122.000000000,89.825,1980.5,2043.0,1616.9,298.90,3477.8,969.57,5.5488,5952.6,2708.5,3360.8,2032.1,0.0000,-6646.5,-6902.2,-1387.9,-2185.0,-2217.2,-15896.,-113.38,-19530.,-6218.0,-4132.4,-2491.7,87.113,2377.2,2180.0,1692.8,348.40,3707.8,1686.6,55.026,7065.3,4476.2,4282.2,3691.3,0.0000,-364.94,-112.82,-91.222,-43.929,-113.27,-587.69,-2.5128,-1064.7,-1545.2,-749.87,-1223.5
1123.000000000,89.963,1983.5,2045.0,1611.5,299.35,3464.4,969.56,5.5494,5942.6,2708.7,3360.7,2032.3,0.0000,-6644.1,-6900.9,-1385.9,-2184.2,-2213.8,-15894.,-113.33,-19528.,-6217.6,-4131.8,-2491.0,65.725,2341.4,2135.0,1671.8,330.31,3675.4,1686.6,0.0000,7032.4,4449.7,4252.8,3658.0,0.0000,-364.83,-111.84,-91.007,-43.817,-112.60,-587.69,0.0000,-1064.3,-1545.1,-749.70,-1222.7
1124.000000000,89.965,1984.0,2045.9,1607.4,299.28,3451.6,969.57,5.5499,5933.6,2709.0,3360.7,2032.4,0.0000,-6641.8,-6899.9,-1383.9,-2183.4,-2210.5,-15892.,-113.28,-19526.,-6217.2,-4131.3,-2490.2,65.649,2338.7,2132.5,1664.5,329.83,3657.1,1686.6,0.0000,7021.3,4449.7,4252.8,3658.0,0.0000,-364.37,-111.68,-90.714,-43.766,-111.94,-587.69,0.0000,-1064.1,-1545.1,-749.69,-1222.5
1125.000000000,89.964,1982.8,2044.3,1602.5,299.33,3437.5,969.57,5.5504,5924.2,2709.2,3360.8,2032.5,0.0000,-6639.4,-6898.7,-1382.0,-2182.7,-2207.3,-15890.,-113.23,-19524.,-6216.7,-4130.7,-2489.4,65.538,2334.8,2128.9,1656.7,329.19,3638.1,1686.6,0.0000,7009.8,4449.7,4252.8,3658.0,0.0000,-363.72,-111.47,-90.391,-43.692,-111.26,-587.69,0.0000,-1064.0,-1545.0,-749.67,-1222.4
1126.000000000,89.957,1980.2,2041.8,1597.0,298.94,3426.9,969.57,5.5509,5914.4,2709.1,3360.8,2032.6,0.0000,-6637.0,-6897.5,-1380.0,-2181.9,-2203.9,-15888.,-113.18,-19522.,-6216.3,-4130.2,-2488.7,65.403,2329.9,2124.5,1648.5,328.43,3618.6,1686.6,0.0000,6997.9,4449.7,4252.8,3658.0,0.0000,-362.93,-111.22,-90.043,-43.602,-110.56,-587.69,0.0000,-1063.9,-1544.9,-749.66,-1222.3
1127.000000000,89.853,1976.9,2038.5,1590.6,298.34,3410.7,969.56,5.5514,5905.0,2709.1,3360.8,2032.7,0.0000,-6634.4,-6896.3,-1378.0,-2181.1,-2200.5,-15887.,-113.13,-19519.,-6215.8,-4129.7,-2487.9,65.253,2324.6,2119.7,1640.2,327.60,3598.6,1686.6,0.0000,6985.8,4449.7,4252.8,3658.0,0.0000,-362.06,-110.94,-89.682,-43.502,-109.85,-587.69,0.0000,-1063.8,-1544.8,-749.65,-1222.2
1128.000000000,89.738,1973.0,2034.6,1583.7,297.69,3394.2,969.52,5.5519,5896.1,2709.2,3360.7,2032.7,0.0000,-6631.6,-6894.9,-1375.9,-2180.3,-2197.1,-15885.,-113.08,-19517.,-6215.4,-4129.1,-2487.1,65.101,2319.2,2114.7,1632.0,326.77,3579.0,1686.6,0.0000,6973.9,4449.7,4252.8,3658.0,0.0000,-361.18,-110.66,-89.323,-43.401,-109.15,-587.69,0.0000,-1063.7,-1544.7,-749.63,-1222.0
1129.000000000,89.622,1969.1,2031.0,1576.2,297.00,3379.3,969.52,5.5524,5888.4,2709.2,3360.7,2032.8,0.0000,-6628.7,-6893.5,-1373.8,-2179.5,-2193.7,-15883.,-113.03,-19515.,-6215.0,-4128.6,-2486.4,64.973,2314.6,2110.6,1624.4,326.05,3560.7,1686.6,0.0000,6962.8,4449.7,4252.8,3658.0,0.0000,-360.43,-110.42,-88.996,-43.315,-108.48,-587.69,0.0000,-1063.5,-1544.6,-749.62,-1221.9
1130.000000000,89.482,1966.0,2027.4,1568.5,296.34,3364.8,969.52,5.5529,5879.5,2709.3,3360.7,2032.8,0.0000,-6625.8,-6892.1,-1371.6,-2178.6,-2190.2,-15881.,-112.98,-19513.,-6214.5,-4128.0,-2485.6,64.859,2310.6,2106.8,1617.1,325.40,3543.1,1686.6,0.0000,6952.1,4449.7,4252.8,3658.0,0.0000,-359.75,-110.20,-88.688,-43.239,-107.84,-587.69,0.0000,-1063.4,-1544.5,-749.60,-1221.8
1131.000000000,89.350,1963.0,2023.7,1561.5,295.70,3348.9,969.53,5.5562,5869.9,2709.4,3360.7,2032.8,0.0000,-6622.7,-6890.6,-1369.5,-2177.8,-2186.9,-15879.,-112.93,-19511.,-6214.1,-4127.5,-2484.8,64.737,2306.2,2102.9,1609.8,324.71,3525.4,1686.6,0.0000,6941.4,4449.7,4252.8,3658.0,0.0000,-359.03,-109.97,-88.374,-43.158,-107.19,-587.69,0.0000,-1063.3,-1544.4,-749.59,-1221.7
1132.000000000,89.219,1959.6,2019.9,1554.8,295.09,3332.4,969.51,5.5593,5859.8,2709.6,3360.7,2032.9,0.0000,-6619.6,-6889.1,-1367.3,-2176.9,-2183.5,-15877.,-112.88,-19509.,-6213.7,-4126.9,-2484.1,64.607,2301.6,2098.7,1602.3,323.99,3507.5,1686.6,0.0000,6930.5,4449.7,4252.8,3658.0,0.0000,-358.27,-109.72,-88.052,-43.071,-106.54,-587.69,0.0000,-1063.2,-1544.3,-749.58,-1221.6
1133.000000000,89.090,1956.2,2016.0,1547.8,294.45,3315.6,969.49,5.2356,5849.2,2709.8,3360.6,2033.1,0.0000,-6616.4,-6887.6,-1365.0,-2176.1,-2180.2,-15876.,-112.83,-19507.,-6213.3,-4126.4,-2483.3,64.473,2296.8,2094.3,1594.8,323.25,3489.5,1686.6,0.0000,6919.6,4449.7,4252.8,3658.0,0.0000,-357.48,-109.47,-87.726,-42.982,-105.88,-587.69,0.0000,-1063.1,-1544.2,-749.56,-1221.4
1134.000000000,88.958,1952.4,2011.9,1540.8,293.79,3299.0,969.49,4.6125,5838.6,2709.9,3360.6,2033.2,0.0000,-6613.1,-6886.0,-1362.8,-2175.2,-2177.0,-15874.,-112.78,-19504.,-6212.8,-4125.8,-2482.5,64.331,2291.7,2089.7,1587.2,322.46,3471.4,1686.6,0.0000,6908.6,4449.7,4252.8,3658.0,0.0000,-356.64,-109.20,-87.393,-42.887,-105.22,-587.69,0.0000,-1063.0,-1544.2,-749.55,-1221.3
1135.000000000,88.757,1948.2,2008.0,1533.6,293.10,3282.7,969.49,4.6129,5828.4,2710.0,3360.6,2033.2,0.0000,-6609.7,-6884.5,-1360.5,-2174.4,-2173.9,-15872.,-112.73,-19502.,-6212.4,-4125.2,-2481.8,64.194,2286.9,2085.2,1579.8,321.71,3453.5,1686.6,0.0000,6897.8,4449.7,4252.8,3658.0,0.0000,-355.83,-108.94,-87.067,-42.796,-104.57,-587.69,0.0000,-1062.8,-1544.1,-749.53,-1221.2
1136.000000000,88.605,1944.4,2003.8,1526.5,292.36,3266.5,969.49,4.6132,5818.3,2710.1,3360.6,2033.3,0.0000,-6606.2,-6882.9,-1358.3,-2173.5,-2170.7,-15870.,-112.68,-19500.,-6212.0,-4124.7,-2481.0,64.045,2281.6,2080.4,1572.1,320.89,3435.3,1686.6,0.0000,6886.7,4449.7,4252.8,3658.0,0.0000,-354.96,-108.66,-86.729,-42.697,-103.91,-587.69,0.0000,-1062.7,-1544.0,-749.52,-1221.1
1137.000000000,88.458,1940.1,1999.8,1519.4,291.65,3250.2,969.49,4.6136,5808.1,2710.0,3360.6,2033.3,0.0000,-6602.6,-6881.2,-1356.0,-2172.6,-2167.5,-15868.,-112.63,-19498.,-6211.6,-4124.1,-2480.2,63.886,2275.9,2075.2,1564.3,320.03,3416.7,1686.6,0.0000,6875.5,4449.7,4252.8,3658.0,0.0000,-354.03,-108.36,-86.378,-42.590,-103.21,-587.69,0.0000,-1062.6,-1543.9,-749.50,-1221.0
1138.000000000,88.303,1935.6,1995.3,1512.1,290.93,3237.1,969.49,4.6140,5798.0,2710.3,3360.5,2033.4,0.0000,-6599.0,-6879.5,-1353.7,-2171.7,-2164.3,-15866.,-112.58,-19496.,-6211.1,-4123.6,-2479.5,63.718,2269.9,2069.8,1556.3,319.12,3397.9,1686.6,0.0000,6864.1,4449.7,4252.8,3658.0,0.0000,-353.05,-108.04,-86.019,-42.479,-102.51,-587.69,0.0000,-1062.5,-1543.8,-749.49,-1220.8
1139.000000000,88.141,1931.1,1990.8,1504.9,290.16,3221.9,969.49,4.6144,5788.1,2710.3,3360.5,2033.5,0.0000,-6595.2,-6877.8,-1351.3,-2170.8,-2161.0,-15864.,-112.54,-19493.,-6210.7,-4123.0,-2478.7,63.551,2264.0,2064.4,1548.4,318.22,3379.2,1686.6,0.0000,6852.7,4449.7,4252.8,3658.0,0.0000,-352.07,-107.73,-85.661,-42.367,-101.82,-587.69,0.0000,-1062.4,-1543.7,-749.48,-1220.7
1140.000000000,88.100,1926.2,1986.1,1497.5,289.38,3205.4,969.49,4.6148,5778.1,2710.4,3360.6,2033.6,0.0000,-6591.3,-6876.0,-1349.0,-2169.9,-2157.7,-15862.,-112.49,-19491.,-6210.3,-4122.5,-2477.9,63.382,2258.0,2058.9,1540.5,317.31,3360.5,1686.6,0.0000,6841.4,4449.7,4252.8,3658.0,0.0000,-351.08,-107.41,-85.304,-42.255,-101.12,-587.69,0.0000,-1062.2,-1543.6,-749.46,-1220.6
1141.000000000,87.995,1921.5,1981.0,1490.2,288.59,3188.7,969.49,4.6152,5767.9,2710.4,3360.6,2033.8,0.0000,-6587.3,-6874.2,-1346.6,-2169.0,-2154.3,-15861.,-112.45,-19489.,-6209.9,-4121.9,-2477.2,63.222,2252.2,2053.7,1532.8,316.44,3342.3,1686.6,0.0000,6830.4,4449.7,4252.8,3658.0,0.0000,-350.14,-107.11,-84.958,-42.148,-100.44,-587.69,0.0000,-1062.1,-1543.5,-749.45,-1220.5
1142.000000000,87.859,1916.8,1975.9,1483.0,287.81,3172.1,969.49,4.6156,5757.7,2710.4,3360.6,2033.9,0.0000,-6583.2,-6872.4,-1344.2,-2168.1,-2150.9,-15859.,-112.40,-19486.,-6209.4,-4121.4,-2476.4,63.063,2246.6,2048.5,1525.1,315.58,3324.2,1686.6,0.0000,6819.4,4449.7,4252.8,3658.0,0.0000,-349.20,-106.80,-84.614,-42.042,-99.756,-587.69,0.0000,-1062.0,-1543.4,-749.43,-1220.3
1143.000000000,87.705,1912.0,1971.1,1475.7,286.93,3155.8,969.50,4.6160,5747.7,2710.3,3360.6,2034.0,0.0000,-6579.1,-6870.5,-1341.8,-2167.2,-2147.5,-15857.,-112.35,-19484.,-6209.0,-4120.8,-2475.6,62.896,2240.6,2043.1,1517.3,314.68,3305.9,1686.6,0.0000,6808.3,4449.7,4252.8,3658.0,0.0000,-348.22,-106.49,-84.262,-41.931,-99.068,-587.69,0.0000,-1061.9,-1543.3,-749.42,-1220.2
1144.000000000,87.536,1907.1,1966.3,1468.4,286.14,3139.2,969.50,4.6163,5737.8,2710.1,3360.7,2034.1,0.0000,-6574.8,-6868.6,-1339.4,-2166.2,-2144.0,-15855.,-112.31,-19482.,-6208.6,-4120.2,-2474.9,62.721,2234.4,2037.4,1509.4,313.74,3287.3,1686.6,0.0000,6797.0,4449.7,4252.8,3658.0,0.0000,-347.19,-106.16,-83.901,-41.814,-98.372,-587.69,0.0000,-1061.8,-1543.3,-749.40,-1220.1
1145.000000000,87.364,1902.1,1961.3,1461.1,285.33,3122.6,969.50,4.6167,5727.6,2710.1,3360.7,2034.2,0.0000,-6570.4,-6866.6,-1336.9,-2165.3,-2140.5,-15853.,-112.26,-19479.,-6208.2,-4119.7,-2474.1,62.538,2227.9,2031.5,1501.4,312.76,3268.5,1686.6,0.0000,6785.6,4449.7,4252.8,3658.0,0.0000,-346.12,-105.81,-83.532,-41.692,-97.668,-587.69,0.0000,-1061.6,-1543.2,-749.39,-1220.0
1146.000000000,87.185,1897.0,1956.4,1453.8,284.49,3105.9,969.50,4.6171,5717.4,2710.3,3360.7,2034.3,0.0000,-6566.0,-6864.7,-1334.4,-2164.3,-2136.9,-15851.,-112.22,-19477.,-6207.7,-4119.1,-2473.4,62.349,2221.2,2025.3,1493.3,311.76,3249.6,1686.6,0.0000,6774.1,4449.7,4252.8,3658.0,0.0000,-345.01,-105.46,-83.157,-41.566,-96.960,-587.69,0.0000,-1061.5,-1543.1,-749.38,-1219.9
1147.000000000,87.000,1891.7,1951.0,1446.3,283.62,3089.3,969.50,4.6175,5707.1,2710.4,3360.7,2034.4,0.0000,-6561.4,-6862.6,-1332.0,-2163.4,-2133.3,-15849.,-112.17,-19475.,-6207.3,-4118.6,-2472.6,62.162,2214.5,2019.2,1485.2,310.76,3230.8,1686.6,0.0000,6762.8,4449.7,4252.8,3658.0,0.0000,-343.91,-105.10,-82.785,-41.441,-96.257,-587.69,0.0000,-1061.4,-1543.0,-749.36,-1219.7
1148.000000000,86.775,1886.9,1946.3,1438.9,282.85,3072.7,969.50,4.7991,5696.9,2710.5,3360.8,2034.5,0.0000,-6556.8,-6860.6,-1329.5,-2162.4,-2129.7,-15847.,-112.13,-19472.,-6206.9,-4118.0,-2471.8,62.154,2214.2,2019.0,1481.3,310.66,3220.6,1686.6,0.0000,6756.6,4449.7,4253.4,3658.9,0.0000,-343.81,-105.06,-82.646,-41.436,-95.817,-587.69,0.0000,-1061.3,-1542.9,-749.35,-1219.6
1149.000000000,86.676,1887.8,1947.1,1432.3,283.07,3057.9,969.50,4.8169,5686.9,2710.6,3360.7,2034.7,0.0000,-6552.6,-6858.8,-1327.1,-2161.5,-2126.1,-15845.,-112.08,-19470.,-6206.4,-4117.4,-2471.1,73.310,2245.0,2056.7,1486.2,318.43,3224.6,1686.6,3.6032,6758.6,4451.8,4254.1,3659.9,0.0000,-348.30,-106.65,-83.239,-42.008,-95.793,-587.69,-0.16452,-1061.2,-1542.8,-749.34,-1219.5
1150.000000000,86.859,1896.9,1954.4,1427.3,284.50,3045.4,969.48,4.8174,5677.7,2710.7,3360.8,2034.8,0.0000,-6549.4,-6857.5,-1324.8,-2160.7,-2122.5,-15843.,-112.04,-19468.,-6206.0,-4116.9,-2470.3,63.188,2251.0,2052.6,1481.1,315.40,3208.4,1686.6,0.0000,6748.9,4449.7,4252.8,3658.0,0.0000,-349.42,-106.75,-83.170,-42.125,-95.175,-587.69,0.0000,-1061.1,-1542.7,-749.32,-1219.4
1151.000000000,87.105,1903.5,1960.7,1423.8,285.14,3033.5,969.45,4.8179,5668.9,2710.9,3360.8,2034.9,0.0000,-6546.6,-6856.6,-1322.5,-2159.9,-2119.0,-15841.,-111.99,-19465.,-6205.6,-4116.3,-2469.6,63.219,2252.1,2053.6,1475.0,315.44,3192.3,1686.6,0.0000,6739.1,4449.7,4252.8,3658.0,0.0000,-349.54,-106.78,-82.978,-42.146,-94.554,-587.69,0.0000,-1061.0,-1542.6,-749.30,-1219.2
1152.000000000,87.258,1906.0,1963.3,1419.9,285.88,3020.4,969.44,4.8184,5659.9,2711.2,3360.8,2035.0,0.0000,-6544.0,-6855.7,-1320.2,-2159.2,-2115.5,-15839.,-111.95,-19463.,-6205.2,-4115.7,-2468.8,63.181,2250.8,2052.3,1468.6,315.15,3176.0,1686.6,0.0000,6729.3,4449.7,4252.8,3658.0,0.0000,-349.29,-106.69,-82.739,-42.121,-93.930,-587.69,0.0000,-1060.9,-1542.5,-749.29,-1219.1
1153.000000000,87.499,1906.0,1963.8,1415.3,286.01,3006.5,969.43,4.0993,5650.7,2711.3,3360.8,2035.1,0.0000,-6541.4,-6854.7,-1318.0,-2158.4,-2111.9,-15837.,-111.90,-19460.,-6204.8,-4115.2,-2468.0,63.099,2247.9,2049.7,1461.8,314.66,3159.4,1686.6,0.0000,6719.2,4449.7,4252.8,3658.0,0.0000,-348.79,-106.53,-82.466,-42.066,-93.296,-587.69,0.0000,-1060.8,-1542.5,-749.28,-1219.0
1154.000000000,87.620,1904.7,1962.9,1409.7,285.71,2992.0,969.43,3.8880,5641.8,2711.4,3360.9,2035.1,0.0000,-6538.7,-6853.6,-1315.7,-2157.6,-2108.2,-15835.,-111.86,-19458.,-6204.3,-4114.6,-2467.3,62.979,2243.6,2045.8,1454.7,313.99,3142.3,1686.6,0.0000,6708.8,4449.7,4252.8,3658.0,0.0000,-348.08,-106.31,-82.160,-41.986,-92.646,-587.69,0.0000,-1060.7,-1542.4,-749.26,-1218.9
1155.000000000,87.529,1902.2,1960.1,1404.1,285.19,2977.1,969.43,3.8973,5633.4,2711.5,3360.9,2035.3,0.0000,-6535.8,-6852.5,-1313.5,-2156.7,-2104.6,-15833.,-111.81,-19456.,-6203.9,-4114.1,-2466.5,62.832,2238.4,2041.0,1447.4,313.19,3124.9,1686.6,0.0000,6698.2,4449.7,4252.8,3658.0,0.0000,-347.22,-106.04,-81.834,-41.888,-91.988,-587.69,0.0000,-1060.5,-1542.3,-749.25,-1218.8
1156.000000000,87.581,1898.8,1957.2,1397.6,284.57,2963.2,969.43,3.9137,5626.1,2711.7,3360.9,2035.4,0.0000,-6532.8,-6851.3,-1311.1,-2155.9,-2100.8,-15831.,-111.77,-19453.,-6203.5,-4113.5,-2465.8,62.682,2233.0,2036.1,1440.1,312.38,3107.7,1686.6,0.0000,6687.8,4449.7,4252.8,3658.0,0.0000,-346.35,-105.76,-81.508,-41.788,-91.338,-587.69,0.0000,-1060.4,-1542.2,-749.23,-1218.6
1157.000000000,87.444,1895.3,1953.9,1390.9,283.89,2949.9,969.43,3.9148,5618.5,2711.6,3361.0,2035.5,0.0000,-6529.7,-6850.0,-1308.8,-2155.0,-2097.1,-15829.,-111.72,-19451.,-6203.1,-4112.9,-2465.0,62.531,2227.6,2031.2,1433.0,311.56,3090.9,1686.6,0.0000,6677.6,4449.7,4252.8,3658.0,0.0000,-345.46,-105.48,-81.186,-41.687,-90.698,-587.69,0.0000,-1060.3,-1542.1,-749.22,-1218.5
1158.000000000,87.296,1891.7,1950.4,1384.4,283.17,2936.2,969.43,3.9151,5610.2,2711.6,3361.0,2035.6,0.0000,-6526.4,-6848.6,-1306.4,-2154.2,-2093.3,-15827.,-111.68,-19448.,-6202.7,-4112.4,-2464.3,62.368,2221.8,2025.9,1425.8,310.69,3074.0,1686.6,0.0000,6667.4,4449.7,4252.8,3658.0,0.0000,-344.51,-105.18,-80.855,-41.579,-90.055,-587.69,0.0000,-1060.2,-1542.0,-749.20,-1218.4
1159.000000000,87.137,1887.7,1946.4,1378.3,282.43,2921.4,969.40,3.9118,5601.6,2711.6,3361.1,2035.7,0.0000,-6523.0,-6847.1,-1304.0,-2153.3,-2089.4,-15825.,-111.63,-19446.,-6202.2,-4111.8,-2463.5,62.201,2215.9,2020.5,1418.5,309.80,3057.1,1686.6,0.0000,6657.1,4449.7,4252.8,3658.0,0.0000,-343.54,-104.87,-80.522,-41.468,-89.415,-587.69,0.0000,-1060.1,-1541.9,-749.19,-1218.3
1160.000000000,86.972,1883.8,1942.0,1371.9,281.67,2906.2,969.40,3.8820,5592.5,2711.6,3361.0,2035.8,0.0000,-6519.4,-6845.6,-1301.6,-2152.4,-2085.6,-15823.,-111.59,-19443.,-6201.8,-4111.2,-2462.7,62.034,2209.9,2015.1,1411.4,308.91,3040.4,1686.6,0.0000,6647.1,4449.7,4252.8,3658.0,0.0000,-342.57,-104.56,-80.192,-41.356,-88.781,-587.69,0.0000,-1060.0,-1541.8,-749.17,-1218.2
1161.000000000,86.917,1879.6,1937.6,1365.2,280.89,2890.8,969.40,3.8824,5583.2,2711.7,3361.0,2035.9,0.0000,-6515.7,-6844.1,-1299.2,-2151.5,-2081.7,-15821.,-111.54,-19441.,-6201.4,-4110.7,-2462.0,61.857,2203.6,2009.4,1404.2,307.98,3023.6,1686.6,0.0000,6636.9,4449.7,4252.8,3658.0,0.0000,-341.54,-104.23,-79.853,-41.238,-88.142,-587.69,0.0000,-1059.8,-1541.7,-749.16,-1218.0
1162.000000000,86.816,1875.0,1932.8,1358.5,280.04,2875.6,969.40,3.8828,5573.7,2711.6,3361.0,2036.0,0.0000,-6511.8,-6842.4,-1296.7,-2150.6,-2077.8,-15819.,-111.50,-19438.,-6200.9,-4110.1,-2461.2,61.671,2197.0,2003.3,1396.8,306.99,3006.5,1686.6,0.0000,6626.5,4449.7,4252.8,3658.0,0.0000,-340.45,-103.89,-79.504,-41.114,-87.495,-587.69,0.0000,-1059.7,-1541.7,-749.14,-1217.9
1163.000000000,86.737,1876.9,1934.0,1352.1,280.32,2862.1,969.40,3.8832,5564.6,2711.6,3361.0,2036.1,0.0000,-6508.2,-6841.0,-1294.4,-2149.7,-2073.9,-15817.,-111.45,-19436.,-6200.5,-4109.5,-2460.5,106.72,2250.4,2081.6,1415.6,318.63,3038.7,1686.6,2.6561,6646.4,4452.7,4255.6,3661.2,0.0000,-347.85,-106.87,-80.799,-42.043,-88.274,-587.69,-0.12128,-1059.8,-1541.6,-749.14,-1217.9
1164.000000000,87.698,1896.5,1950.3,1348.5,283.48,2853.6,969.38,3.8836,5556.9,2711.7,3361.1,2036.2,0.0000,-6506.4,-6840.6,-1292.3,-2149.0,-2070.1,-15815.,-111.41,-19434.,-6200.1,-4109.0,-2459.7,391.96,2337.4,2529.4,1433.8,343.19,3068.8,1686.6,0.0000,6661.9,4455.1,4270.2,3675.8,0.0000,-355.30,-117.75,-81.910,-43.051,-88.695,-587.69,0.0000,-1059.9,-1541.5,-749.20,-1218.1
1165.000000000,88.713,1927.9,1979.3,1350.4,287.83,2851.8,969.37,3.8923,5550.7,2711.8,3361.2,2036.3,0.0000,-6506.7,-6841.5,-1290.5,-2148.6,-2066.6,-15813.,-111.37,-19431.,-6199.6,-4108.4,-2459.0,469.92,2641.4,2647.2,1483.8,390.49,3158.8,1686.7,33.201,6717.6,4474.6,4300.2,3706.1,0.0000,-365.99,-122.13,-83.965,-44.533,-90.535,-587.69,-1.5159,-1060.3,-1541.4,-749.34,-1218.6
1166.000000000,90.055,1971.1,2019.3,1358.8,294.94,2862.3,969.37,3.9077,5547.9,2711.9,3361.1,2036.4,0.0000,-6509.7,-6843.9,-1289.3,-2148.4,-2063.7,-15811.,-111.33,-19429.,-6199.2,-4107.8,-2458.2,745.17,2966.7,2876.7,1597.5,462.50,3381.1,1687.9,332.13,6858.8,4510.3,4347.5,3752.9,0.0000,-379.42,-129.40,-87.802,-46.475,-95.781,-587.71,-15.165,-1061.5,-1541.3,-749.57,-1219.5
1167.000000000,92.070,2021.5,2066.8,1380.4,303.26,2892.0,969.37,3.9106,5551.0,2712.0,3361.2,2036.4,0.0000,-6515.7,-6847.8,-1288.8,-2148.5,-2061.4,-15809.,-111.29,-19426.,-6198.8,-4107.3,-2457.5,518.86,2752.1,2645.9,1663.3,518.63,3511.1,1702.0,160.58,6934.7,4562.6,4402.2,3804.5,0.0000,-388.10,-126.17,-89.806,-47.867,-98.017,-587.92,-7.3320,-1062.2,-1541.2,-749.83,-1220.4
1168.000000000,93.846,2066.2,2111.1,1410.0,311.17,2931.2,969.37,3.9111,5558.5,2712.1,3361.6,2036.6,0.0000,-6523.6,-6852.7,-1288.8,-2148.7,-2060.1,-15807.,-111.25,-19424.,-6198.4,-4106.7,-2456.7,71.400,2543.6,2319.3,1602.5,370.64,3429.7,1686.6,0.0000,6878.4,4451.6,4260.7,3663.6,0.0000,-394.22,-120.43,-91.382,-47.696,-99.066,-587.69,0.0000,-1061.0,-1541.1,-749.10,-1217.3
1169.000000000,95.443,2098.2,2143.4,1439.5,316.96,2968.2,969.37,3.9115,5568.9,2712.3,3361.5,2036.8,0.0000,-6532.4,-6857.8,-1289.4,-2149.0,-2059.3,-15805.,-111.21,-19422.,-6197.9,-4106.1,-2456.0,71.557,2549.2,2324.4,1620.6,365.14,3476.4,1686.6,0.0000,6908.1,4450.5,4256.8,3660.6,0.0000,-395.17,-120.77,-92.168,-47.760,-100.50,-587.69,0.0000,-1061.1,-1541.1,-749.06,-1217.2
1170.000000000,96.352,2113.7,2162.1,1468.9,319.81,3002.5,969.37,3.9162,5580.4,2712.4,3361.8,2037.0,0.0000,-6540.8,-6862.5,-1290.2,-2149.2,-2058.6,-15803.,-111.16,-19420.,-6197.5,-4105.6,-2455.2,71.479,2546.4,2321.9,1636.3,358.51,3518.2,1686.6,0.0000,6935.1,4449.7,4253.5,3658.4,0.0000,-394.84,-120.72,-92.728,-47.668,-101.79,-587.69,0.0000,-1061.3,-1541.0,-749.03,-1217.0
1171.000000000,96.786,2120.4,2172.5,1492.7,321.11,3037.2,969.37,3.9141,5597.5,2712.5,3362.0,2037.2,0.0000,-6548.5,-6866.6,-1291.3,-2149.2,-2058.0,-15801.,-111.12,-19418.,-6197.1,-4105.0,-2454.5,71.309,2540.3,2316.4,1651.4,355.88,3559.3,1686.6,0.0000,6960.6,4449.7,4252.8,3658.0,0.0000,-393.99,-120.50,-93.172,-47.541,-102.98,-587.69,0.0000,-1061.4,-1540.9,-749.01,-1216.9
1172.000000000,96.834,2123.0,2177.3,1514.5,321.05,3070.7,969.37,3.9145,5619.4,2712.4,3362.0,2037.4,0.0000,-6555.3,-6870.0,-1292.6,-2149.1,-2057.4,-15799.,-111.08,-19416.,-6196.6,-4104.4,-2453.7,71.101,2532.9,2309.6,1665.5,354.88,3598.4,1686.6,0.0000,6984.5,4449.7,4252.8,3658.0,0.0000,-392.93,-120.21,-93.551,-47.401,-104.09,-587.69,0.0000,-1061.5,-1540.8,-749.00,-1216.8
1173.000000000,96.648,2122.4,2179.2,1532.3,320.58,3110.4,969.38,3.9149,5651.9,2712.5,3362.0,2037.6,0.0000,-6561.4,-6872.9,-1293.9,-2148.9,-2056.9,-15797.,-111.03,-19414.,-6196.2,-4103.9,-2453.0,70.837,2523.5,2301.1,1677.5,353.87,3632.5,1686.6,0.0000,7005.3,4449.7,4252.8,3658.0,0.0000,-391.55,-119.82,-93.826,-47.225,-105.06,-587.69,0.0000,-1061.6,-1540.7,-748.98,-1216.7
1174.000000000,96.497,2123.0,2180.3,1548.6,320.23,3158.2,969.38,3.9153,5687.2,2712.5,3362.2,2037.7,0.0000,-6566.8,-6875.3,-1295.1,-2148.7,-2056.5,-15795.,-110.99,-19412.,-6195.8,-4103.3,-2452.2,70.971,2675.1,2464.1,1813.8,502.15,3837.1,1686.6,198.52,7149.6,4561.2,4398.6,3796.4,0.0000,-392.61,-123.48,-94.661,-48.222,-107.39,-587.69,-9.0644,-1063.3,-1540.6,-749.71,-1219.4
1175.000000000,96.546,2125.4,2181.6,1565.3,320.30,3208.8,969.37,3.9156,5719.2,2712.4,3362.4,2037.9,0.0000,-6571.8,-6877.6,-1296.4,-2148.4,-2056.2,-15793.,-110.94,-19410.,-6195.4,-4102.7,-2451.5,70.836,2523.5,2301.0,1711.9,354.46,3721.7,1686.6,0.0000,7059.5,4449.7,4252.8,3658.0,0.0000,-391.70,-119.92,-95.001,-47.224,-107.63,-587.69,0.0000,-1061.8,-1540.6,-748.95,-1216.4
1176.000000000,96.755,2125.7,2181.0,1583.2,320.03,3250.9,969.37,3.9160,5747.9,2712.5,3362.6,2038.0,0.0000,-6576.2,-6879.7,-1297.7,-2148.1,-2056.0,-15791.,-110.90,-19409.,-6194.9,-4102.2,-2450.8,70.644,2516.7,2294.8,1721.8,353.75,3749.8,1686.6,0.0000,7076.6,4449.7,4252.8,3658.0,0.0000,-390.70,-119.64,-95.244,-47.096,-108.44,-587.69,0.0000,-1061.9,-1540.5,-748.94,-1216.3
1177.000000000,96.484,2124.2,2178.7,1599.0,319.71,3285.9,969.37,3.9164,5771.8,2712.6,3362.9,2038.1,0.0000,-6579.8,-6881.5,-1299.0,-2147.8,-2055.9,-15789.,-110.86,-19407.,-6194.5,-4101.6,-2450.0,70.414,2508.5,2287.3,1730.1,352.83,3773.9,1686.6,0.0000,7091.3,4449.7,4252.8,3658.0,0.0000,-389.49,-119.28,-95.410,-46.943,-109.13,-587.69,0.0000,-1061.9,-1540.4,-748.93,-1216.2
1178.000000000,96.312,2120.4,2175.7,1611.8,319.00,3315.6,969.37,3.9168,5792.2,2712.9,3363.3,2038.3,0.0000,-6582.8,-6883.0,-1300.2,-2147.4,-2055.9,-15787.,-110.81,-19406.,-6194.1,-4101.0,-2449.3,70.139,2498.7,2278.4,1736.6,351.68,3793.8,1686.6,0.0000,7103.5,4449.7,4252.8,3658.0,0.0000,-388.02,-118.85,-95.490,-46.760,-109.70,-587.69,0.0000,-1062.0,-1540.3,-748.91,-1216.1
1179.000000000,96.072,2115.0,2171.9,1622.0,318.17,3342.8,969.37,3.9172,5810.8,2713.0,3363.2,2038.5,0.0000,-6585.2,-6884.2,-1301.5,-2147.0,-2055.8,-15785.,-110.77,-19404.,-6193.7,-4100.5,-2448.5,69.882,2489.5,2270.0,1742.5,350.60,3812.1,1686.6,0.0000,7114.7,4449.7,4252.8,3658.0,0.0000,-386.64,-118.44,-95.561,-46.588,-110.23,-587.69,0.0000,-1062.0,-1540.2,-748.90,-1216.0
1180.000000000,95.822,2109.4,2167.4,1630.6,317.42,3369.4,969.37,3.9175,5829.0,2713.1,3363.2,2038.7,0.0000,-6587.2,-6885.3,-1302.6,-2146.6,-2055.8,-15783.,-110.72,-19403.,-6193.2,-4099.9,-2447.8,69.626,2480.4,2261.7,1747.5,349.51,3828.1,1686.6,0.0000,7124.5,4449.7,4252.8,3658.0,0.0000,-385.26,-118.02,-95.602,-46.417,-110.69,-587.69,0.0000,-1062.0,-1540.1,-748.88,-1215.9
1181.000000000,95.560,2103.5,2162.8,1637.7,316.45,3396.4,969.34,3.9179,5848.4,2713.1,3363.2,2038.8,0.0000,-6588.8,-6886.0,-1303.7,-2146.1,-2055.9,-15781.,-110.68,-19402.,-6192.8,-4099.4,-2447.0,69.356,2470.8,2252.9,1751.5,348.34,3841.3,1686.6,0.0000,7132.6,4449.7,4252.8,3658.0,0.0000,-383.81,-117.58,-95.598,-46.238,-111.06,-587.69,0.0000,-1062.1,-1540.0,-748.87,-1215.7
1182.000000000,95.291,2097.1,2156.4,1644.6,315.46,3421.1,969.34,3.9183,5864.2,2713.6,3363.1,2039.1,0.0000,-6589.9,-6886.5,-1304.7,-2145.6,-2056.0,-15779.,-110.64,-19400.,-6192.4,-4098.8,-2446.3,69.062,2460.3,2243.4,1754.0,347.04,3851.3,1686.6,0.0000,7138.7,4449.7,4252.8,3658.0,0.0000,-382.20,-117.10,-95.535,-46.041,-111.35,-587.69,0.0000,-1062.1,-1540.0,-748.85,-1215.6
1183.000000000,94.779,2089.7,2148.6,1650.9,314.44,3441.0,969.33,3.9186,5877.3,2713.9,3363.4,2039.2,0.0000,-6590.5,-6886.7,-1305.5,-2145.1,-2056.1,-15777.,-110.59,-19399.,-6192.0,-4098.2,-2445.5,68.789,2450.6,2234.5,1756.2,345.82,3860.2,1686.6,0.0000,7144.1,4449.7,4252.8,3658.0,0.0000,-380.71,-116.64,-95.470,-45.859,-111.60,-587.69,0.0000,-1062.1,-1539.9,-748.84,-1215.5
1184.000000000,94.468,2082.1,2140.7,1655.9,313.51,3457.1,969.30,3.9190,5889.6,2714.1,3363.2,2039.4,0.0000,-6590.5,-6886.7,-1306.3,-2144.5,-2056.2,-15776.,-110.55,-19398.,-6191.6,-4097.7,-2444.8,68.509,2440.6,2225.4,1757.6,344.56,3866.8,1686.6,0.0000,7148.3,4449.7,4252.8,3658.0,0.0000,-379.18,-116.17,-95.374,-45.673,-111.78,-587.69,0.0000,-1062.1,-1539.8,-748.83,-1215.4
1185.000000000,93.947,2074.3,2132.7,1660.0,312.41,3470.0,969.30,3.2377,5900.9,2714.5,3362.7,2039.5,0.0000,-6590.1,-6886.3,-1307.0,-2143.9,-2056.4,-15774.,-110.50,-19397.,-6191.2,-4097.1,-2444.0,68.203,2429.7,2215.5,1757.6,343.15,3870.4,1686.6,0.0000,7150.5,4449.7,4252.8,3658.0,0.0000,-377.49,-115.65,-95.217,-45.468,-111.88,-587.69,0.0000,-1062.0,-1539.7,-748.81,-1215.3
1186.000000000,93.612,2066.3,2124.0,1663.0,311.25,3482.5,969.30,2.9672,5910.1,2714.3,3362.6,2039.6,0.0000,-6589.3,-6885.8,-1307.6,-2143.2,-2056.5,-15772.,-110.46,-19396.,-6190.7,-4096.6,-2443.3,67.886,2418.4,2205.2,1756.7,341.68,3871.6,1686.6,0.0000,7151.3,4449.7,4252.8,3658.0,0.0000,-375.73,-115.10,-95.024,-45.257,-111.90,-587.69,0.0000,-1062.0,-1539.6,-748.80,-1215.2
1187.000000000,93.307,2058.0,2115.6,1665.1,310.08,3492.5,969.30,2.9675,5918.5,2714.4,3362.7,2039.4,0.0000,-6588.0,-6885.0,-1308.1,-2142.6,-2056.7,-15770.,-110.42,-19395.,-6190.3,-4096.0,-2442.6,67.603,2408.3,2196.0,1755.7,340.37,3872.2,1686.6,0.0000,7151.7,4449.7,4252.8,3658.0,0.0000,-374.17,-114.61,-94.845,-45.069,-111.91,-587.69,0.0000,-1062.0,-1539.5,-748.79,-1215.1
1188.000000000,93.013,2050.0,2109.6,1666.2,308.87,3501.0,969.30,2.9678,5925.8,2714.1,3362.7,2039.6,0.0000,-6586.5,-6884.0,-1308.5,-2141.9,-2056.9,-15768.,-110.37,-19394.,-6189.9,-4095.5,-2441.8,67.368,2399.9,2188.4,1755.4,339.28,3873.9,1686.6,0.0000,7152.8,4449.7,4252.8,3658.0,0.0000,-372.85,-114.20,-94.711,-44.912,-111.94,-587.69,0.0000,-1062.0,-1539.5,-748.77,-1214.9
1189.000000000,92.835,2042.9,2104.8,1666.6,307.77,3509.3,969.30,2.9682,5932.6,2714.9,3362.4,2039.7,0.0000,-6584.7,-6882.8,-1308.8,-2141.1,-2057.0,-15766.,-110.33,-19393.,-6189.5,-4094.9,-2441.1,67.121,2391.1,2180.3,1754.2,338.13,3873.6,1686.6,0.0000,7152.7,4449.7,4252.8,3658.0,0.0000,-371.47,-113.77,-94.543,-44.747,-111.92,-587.69,0.0000,-1061.9,-1539.4,-748.76,-1214.8
1190.000000000,92.603,2036.3,2099.3,1666.5,306.75,3515.1,969.28,2.9685,5940.4,2715.5,3362.2,2040.1,0.0000,-6582.9,-6881.5,-1309.1,-2140.4,-2057.2,-15765.,-110.28,-19391.,-6189.2,-4094.4,-2440.3,66.860,2381.8,2171.8,1752.2,336.90,3871.3,1686.6,0.0000,7151.3,4449.7,4252.8,3658.0,0.0000,-370.00,-113.30,-94.340,-44.573,-111.83,-587.69,0.0000,-1061.9,-1539.3,-748.74,-1214.7
1191.000000000,92.603,2028.8,2092.0,1666.1,305.71,3519.0,969.27,2.9688,5947.4,2715.2,3362.1,2040.2,0.0000,-6580.8,-6880.1,-1309.2,-2139.6,-2057.2,-15763.,-110.24,-19390.,-6188.8,-4093.8,-2439.6,66.576,2371.7,2162.6,1749.1,335.54,3866.6,1686.6,0.0000,7148.5,4449.7,4252.8,3658.0,0.0000,-368.41,-112.80,-94.090,-44.384,-111.67,-587.69,0.0000,-1061.8,-1539.2,-748.73,-1214.6
1192.000000000,92.541,2020.9,2085.1,1665.5,304.59,3523.2,969.27,2.9691,5951.5,2715.0,3361.9,2040.1,0.0000,-6578.5,-6878.5,-1309.3,-2138.9,-2057.2,-15761.,-110.20,-19389.,-6188.4,-4093.3,-2438.9,66.284,2361.3,2153.1,1745.4,334.13,3860.1,1686.6,0.0000,7144.6,4449.7,4252.8,3658.0,0.0000,-366.76,-112.28,-93.811,-44.189,-111.46,-587.69,0.0000,-1061.8,-1539.1,-748.71,-1214.5
1193.000000000,92.259,2012.7,2078.7,1664.1,303.44,3525.0,969.27,2.9694,5955.6,2715.0,3362.0,2040.1,0.0000,-6576.0,-6876.7,-1309.2,-2138.0,-2057.3,-15760.,-110.15,-19388.,-6188.0,-4092.7,-2438.1,66.012,2351.6,2144.3,1741.6,332.82,3853.4,1686.6,0.0000,7140.6,4449.7,4252.8,3658.0,0.0000,-365.23,-111.79,-93.543,-44.008,-111.24,-587.69,0.0000,-1061.7,-1539.0,-748.70,-1214.4
1194.000000000,91.981,2004.5,2071.4,1661.8,302.29,3525.8,969.27,2.9697,5957.6,2715.0,3362.1,2040.4,0.0000,-6573.3,-6874.7,-1309.1,-2137.2,-2057.4,-15758.,-110.11,-19387.,-6187.6,-4092.2,-2437.4,65.731,2341.6,2135.2,1737.2,331.46,3845.2,1686.6,0.0000,7135.6,4449.7,4252.8,3658.0,0.0000,-363.63,-111.29,-93.248,-43.821,-110.98,-587.69,0.0000,-1061.7,-1539.0,-748.69,-1214.2
1195.000000000,91.696,1996.1,2063.4,1658.7,301.11,3524.8,969.27,3.0163,5958.6,2715.0,3362.0,2040.4,0.0000,-6570.3,-6872.7,-1308.9,-2136.4,-2057.4,-15756.,-110.06,-19386.,-6187.2,-4091.6,-2436.6,65.448,2331.6,2126.0,1732.3,330.08,3835.8,1686.6,0.0000,7130.0,4449.7,4252.8,3658.0,0.0000,-362.03,-110.78,-92.936,-43.632,-110.67,-587.69,0.0000,-1061.6,-1538.9,-748.67,-1214.1
1196.000000000,91.411,1987.8,2055.6,1655.2,299.95,3524.2,969.27,4.7498,5959.1,2715.1,3362.0,2040.5,0.0000,-6566.9,-6870.7,-1308.5,-2135.5,-2057.3,-15755.,-110.02,-19385.,-6186.8,-4091.1,-2435.9,65.174,2321.8,2117.1,1727.3,328.73,3825.7,1686.6,0.0000,7123.9,4449.7,4252.8,3658.0,0.0000,-360.47,-110.28,-92.622,-43.450,-110.34,-587.69,0.0000,-1061.5,-1538.8,-748.66,-1214.0
1197.000000000,91.131,1979.4,2048.0,1651.2,298.78,3521.0,969.28,4.8410,5958.2,2715.2,3362.0,2040.6,0.0000,-6563.4,-6868.6,-1308.1,-2134.6,-2057.1,-15753.,-109.98,-19384.,-6186.4,-4090.5,-2435.2,64.896,2311.9,2108.0,1721.7,327.36,3814.4,1686.6,0.0000,7117.1,4449.7,4252.8,3658.0,0.0000,-358.88,-109.78,-92.289,-43.264,-109.99,-587.69,0.0000,-1061.5,-1538.7,-748.64,-1213.9
1198.000000000,90.849,1971.1,2039.8,1646.9,297.58,3518.2,969.28,3.4436,5956.3,2715.3,3362.1,2040.7,0.0000,-6559.6,-6866.4,-1307.6,-2133.7,-2056.8,-15751.,-109.93,-19382.,-6186.0,-4089.9,-2434.4,64.597,2301.2,2098.3,1715.4,325.88,3801.3,1686.6,0.0000,7109.2,4449.7,4252.8,3658.0,0.0000,-357.18,-109.24,-91.919,-43.064,-109.58,-587.69,0.0000,-1061.4,-1538.6,-748.63,-1213.8
1199.000000000,90.558,1966.8,2034.9,1642.5,297.01,3513.4,969.28,3.4439,5953.8,2715.4,3362.0,2040.8,0.0000,-6555.8,-6864.3,-1307.1,-2132.9,-2056.4,-15749.,-109.89,-19381.,-6185.6,-4089.4,-2433.7,91.126,2327.1,2131.9,1719.0,336.30,3804.3,1686.6,0.0000,7110.9,4449.7,4252.8,3658.0,0.0000,-360.28,-110.49,-92.334,-43.491,-109.63,-587.69,0.0000,-1061.4,-1538.5,-748.61,-1213.7
1200.000000000,90.688,1969.5,2036.0,1638.7,297.59,3510.6,969.28,2.9465,5951.1,2715.5,3361.8,2040.9,0.0000,-6552.6,-6862.5,-1306.5,-2132.0,-2055.9,-15748.,-109.85,-19380.,-6185.2,-4088.8,-2432.9,65.147,2320.8,2116.2,1713.9,328.38,3791.2,1686.6,0.0000,7103.0,4449.7,4252.8,3658.0,0.0000,-360.12,-110.10,-92.150,-43.431,-109.22,-587.69,0.0000,-1061.3,-1538.4,-748.60,-1213.5
1201.000000000,90.523,1969.6,2036.7,1635.7,297.31,3506.2,969.28,2.5010,5949.7,2715.6,3361.7,2041.0,0.0000,-6549.5,-6861.0,-1305.9,-2131.3,-2055.4,-15746.,-109.81,-19379.,-6184.7,-4088.3,-2432.2,65.010,2315.9,2111.8,1707.7,327.64,3776.8,1686.6,0.0000,7094.2,4449.7,4252.8,3658.0,0.0000,-359.32,-109.84,-91.869,-43.340,-108.76,-587.69,0.0000,-1061.2,-1538.4,-748.58,-1213.4
1202.000000000,90.444,1966.8,2033.8,1632.1,297.31,3499.9,969.28,3.1202,5946.4,2715.6,3361.7,2041.1,0.0000,-6546.5,-6859.3,-1305.3,-2130.5,-2054.8,-15744.,-109.76,-19378.,-6184.3,-4087.8,-2431.5,64.822,2309.2,2105.7,1701.1,326.67,3761.7,1686.6,0.0000,7085.0,4449.7,4252.8,3658.0,0.0000,-358.23,-109.50,-91.545,-43.215,-108.28,-587.69,0.0000,-1061.1,-1538.3,-748.57,-1213.3
1203.000000000,90.516,1983.3,2049.6,1629.5,300.42,3499.6,969.28,3.1875,5943.6,2715.6,3361.6,2041.2,0.0000,-6545.0,-6858.6,-1304.9,-2129.8,-2054.3,-15743.,-109.72,-19377.,-6183.9,-4087.2,-2430.8,434.87,2559.8,2455.0,1779.7,365.23,3908.2,1690.8,51.780,7174.7,4455.3,4259.5,3664.4,0.0000,-382.43,-121.29,-96.268,-46.224,-112.37,-587.75,-2.3642,-1061.7,-1538.2,-748.59,-1213.3
1204.000000000,92.771,2039.7,2096.7,1638.3,309.48,3519.8,969.27,3.1878,5946.3,2715.7,3361.6,2041.3,0.0000,-6547.7,-6860.2,-1305.2,-2129.6,-2054.2,-15741.,-109.69,-19376.,-6183.5,-4086.7,-2430.0,238.89,2882.1,2741.1,1865.3,446.67,4079.0,1708.4,210.16,7296.7,4538.2,4357.2,3774.0,0.0000,-390.27,-128.75,-98.590,-47.573,-115.84,-588.01,-9.5958,-1062.8,-1538.1,-749.07,-1215.4
1205.000000000,94.045,2083.8,2141.6,1663.0,314.95,3555.8,969.24,3.1881,5955.0,2715.7,3361.5,2041.4,0.0000,-6552.7,-6863.4,-1306.0,-2129.7,-2055.0,-15740.,-109.65,-19375.,-6183.1,-4086.1,-2429.3,71.445,2545.2,2320.8,1866.1,482.11,4091.4,1686.6,0.0000,7296.6,4488.5,4289.5,3684.5,0.0000,-394.88,-120.76,-99.584,-48.387,-116.59,-587.69,0.0000,-1062.7,-1538.0,-748.71,-1213.5
1206.000000000,95.484,2110.6,2168.9,1688.0,321.83,3588.9,969.24,3.1884,5965.2,2715.7,3361.5,2041.4,0.0000,-6558.6,-6866.8,-1307.2,-2129.8,-2056.3,-15738.,-109.61,-19374.,-6182.7,-4085.6,-2428.6,71.516,2547.7,2323.1,1854.5,375.17,4074.3,1686.6,0.0000,7280.1,4462.5,4264.6,3665.8,0.0000,-395.32,-120.93,-99.889,-47.772,-117.01,-587.69,0.0000,-1062.3,-1538.0,-748.57,-1213.0
1207.000000000,96.568,2122.0,2184.5,1708.0,324.08,3613.4,969.24,3.1887,5974.7,2715.7,3361.5,2041.6,0.0000,-6564.4,-6869.8,-1308.5,-2129.7,-2057.5,-15736.,-109.57,-19374.,-6182.3,-4085.0,-2427.9,71.367,2542.4,2318.3,1851.9,363.19,4077.6,1686.6,0.0000,7277.3,4452.0,4254.8,3658.9,0.0000,-394.55,-120.72,-99.997,-47.602,-117.42,-587.69,0.0000,-1062.2,-1537.9,-748.51,-1212.8
1208.000000000,96.858,2125.5,2188.8,1722.6,324.72,3630.8,969.24,3.1889,5985.8,2715.8,3361.6,2041.6,0.0000,-6569.4,-6872.3,-1310.0,-2129.6,-2058.4,-15735.,-109.52,-19373.,-6181.9,-4084.5,-2427.1,71.161,2535.1,2311.6,1854.3,358.71,4087.7,1686.6,0.0000,7282.2,4449.7,4252.8,3658.0,0.0000,-393.46,-120.41,-100.04,-47.443,-117.82,-587.69,0.0000,-1062.1,-1537.8,-748.48,-1212.6
1209.000000000,96.833,2124.6,2188.5,1733.6,324.23,3646.1,969.24,3.1892,6004.2,2715.8,3361.6,2041.8,0.0000,-6573.4,-6874.2,-1311.5,-2129.3,-2059.3,-15733.,-109.48,-19372.,-6181.5,-4083.9,-2426.4,70.889,2525.4,2302.7,1856.9,357.18,4098.1,1686.6,0.0000,7288.4,4449.7,4252.8,3658.0,0.0000,-392.01,-119.99,-99.998,-47.259,-118.15,-587.69,0.0000,-1062.1,-1537.7,-748.47,-1212.5
1210.000000000,96.625,2121.1,2187.3,1739.3,323.26,3671.4,969.23,3.1895,6030.8,2715.9,3361.7,2041.9,0.0000,-6576.8,-6875.5,-1312.7,-2129.0,-2060.0,-15731.,-109.44,-19371.,-6181.1,-4083.4,-2425.7,70.618,2515.7,2293.9,1859.5,355.99,4107.7,1686.6,0.0000,7294.3,4449.7,4252.8,3658.0,0.0000,-390.55,-119.56,-99.945,-47.079,-118.45,-587.69,0.0000,-1062.2,-1537.6,-748.45,-1212.4
1211.000000000,96.339,2120.0,2186.1,1742.8,322.24,3702.4,969.21,3.1897,6053.6,2716.0,3361.8,2042.0,0.0000,-6579.7,-6876.4,-1313.7,-2128.6,-2060.7,-15730.,-109.40,-19370.,-6180.7,-4082.9,-2424.9,70.291,2504.1,2283.3,1860.1,354.49,4113.2,1686.6,0.0000,7297.7,4449.7,4252.8,3658.0,0.0000,-388.78,-119.03,-99.800,-46.860,-118.63,-587.69,0.0000,-1062.2,-1537.5,-748.44,-1212.3
1212.000000000,95.966,2114.4,2180.2,1749.5,321.02,3722.9,969.21,3.1900,6070.0,2716.4,3361.8,2042.2,0.0000,-6581.8,-6877.0,-1314.5,-2128.1,-2061.3,-15728.,-109.35,-19369.,-6180.3,-4082.3,-2424.2,69.934,2491.4,2271.7,1859.5,352.85,4115.6,1686.6,0.0000,7299.2,4449.7,4252.8,3658.0,0.0000,-386.84,-118.45,-99.596,-46.623,-118.71,-587.69,0.0000,-1062.1,-1537.5,-748.42,-1212.2
1213.000000000,95.647,2109.5,2173.9,1755.9,320.12,3734.3,969.21,3.1903,6080.5,2716.3,3361.9,2042.4,0.0000,-6583.3,-6877.3,-1315.3,-2127.6,-2061.8,-15726.,-109.31,-19368.,-6179.8,-4081.8,-2423.5,268.35,2496.6,2477.7,1867.2,477.44,4133.8,1686.6,0.0000,7310.2,4449.7,4252.8,3658.0,0.0000,-387.69,-123.00,-99.934,-47.485,-119.26,-587.69,0.0000,-1062.2,-1537.4,-748.41,-1212.1
1214.000000000,95.694,2110.6,2171.2,1759.9,319.69,3743.0,969.21,3.1905,6087.3,2716.4,3361.9,2042.5,0.0000,-6584.5,-6877.7,-1316.1,-2127.1,-2062.3,-15725.,-109.27,-19368.,-6179.4,-4081.2,-2422.8,69.855,2488.5,2269.1,1866.2,352.59,4133.7,1686.6,0.0000,7310.3,4449.7,4252.8,3658.0,0.0000,-386.45,-118.34,-99.782,-46.570,-119.28,-587.69,0.0000,-1062.2,-1537.3,-748.39,-1212.0
1215.000000000,95.473,2107.0,2168.8,1762.4,318.81,3751.2,969.21,3.1908,6092.6,2716.5,3361.9,2042.6,0.0000,-6585.2,-6878.0,-1316.7,-2126.6,-2062.8,-15723.,-109.23,-19367.,-6179.0,-4080.7,-2422.0,69.571,2478.4,2259.9,1864.1,351.26,4131.7,1686.6,0.0000,7309.1,4449.7,4252.8,3658.0,0.0000,-384.90,-117.87,-99.567,-46.380,-119.23,-587.69,0.0000,-1062.1,-1537.2,-748.38,-1211.9
1216.000000000,95.280,2100.9,2163.2,1763.8,318.10,3759.0,969.21,3.1911,6098.8,2716.2,3361.9,2042.7,0.0000,-6585.4,-6878.0,-1317.3,-2126.0,-2063.2,-15722.,-109.18,-19366.,-6178.6,-4080.2,-2421.3,69.267,2467.6,2250.1,1861.6,349.82,4128.5,1686.6,0.0000,7307.2,4449.7,4252.8,3658.0,0.0000,-383.23,-117.36,-99.325,-46.178,-119.15,-587.69,0.0000,-1062.1,-1537.1,-748.36,-1211.8
1217.000000000,95.043,2094.3,2157.3,1765.4,316.99,3765.6,969.22,3.1913,6103.2,2716.2,3361.7,2043.0,0.0000,-6585.2,-6877.9,-1317.8,-2125.4,-2063.7,-15720.,-109.14,-19365.,-6178.2,-4079.6,-2420.6,68.973,2457.1,2240.5,1858.8,348.42,4124.5,1686.6,0.0000,7304.8,4449.7,4252.8,3658.0,0.0000,-381.60,-116.86,-99.076,-45.982,-119.05,-587.69,0.0000,-1062.1,-1537.0,-748.35,-1211.6
1218.000000000,94.715,2086.7,2151.4,1765.8,315.81,3768.5,969.19,3.1916,6105.3,2716.4,3361.6,2043.2,0.0000,-6584.7,-6877.5,-1318.2,-2124.8,-2064.0,-15719.,-109.10,-19364.,-6177.7,-4079.1,-2419.9,68.697,2447.3,2231.5,1856.0,347.11,4120.4,1686.6,0.0000,7302.4,4449.7,4252.8,3658.0,0.0000,-380.08,-116.39,-98.840,-45.798,-118.94,-587.69,0.0000,-1062.1,-1537.0,-748.34,-1211.5
1219.000000000,94.444,2080.5,2143.8,1764.6,314.66,3769.6,969.18,3.1919,6108.7,2716.6,3361.8,2043.4,0.0000,-6583.9,-6877.0,-1318.4,-2124.2,-2064.3,-15717.,-109.06,-19363.,-6177.3,-4078.6,-2419.1,68.438,2438.1,2223.1,1853.2,345.87,4116.0,1686.6,0.0000,7299.7,4449.7,4252.8,3658.0,0.0000,-378.64,-115.94,-98.610,-45.625,-118.82,-587.69,0.0000,-1062.0,-1536.9,-748.32,-1211.4
1220.000000000,94.189,2073.1,2135.9,1762.7,313.52,3771.1,969.18,3.1921,6111.4,2716.5,3361.8,2043.5,0.0000,-6582.6,-6876.3,-1318.6,-2123.5,-2064.5,-15715.,-109.01,-19363.,-6176.9,-4078.0,-2418.4,68.153,2427.9,2213.8,1849.3,344.49,4109.2,1686.6,0.0000,7295.7,4449.7,4252.8,3658.0,0.0000,-377.05,-115.45,-98.331,-45.435,-118.62,-587.69,0.0000,-1062.0,-1536.8,-748.31,-1211.3
1221.000000000,93.905,2065.2,2127.9,1760.7,312.28,3771.5,969.18,3.1924,6112.7,2716.5,3361.8,2043.6,0.0000,-6581.0,-6875.4,-1318.7,-2122.8,-2064.8,-15714.,-108.97,-19362.,-6176.5,-4077.5,-2417.7,67.853,2417.2,2204.1,1844.7,343.04,4100.5,1686.6,0.0000,7290.5,4449.7,4252.8,3658.0,0.0000,-375.38,-114.93,-98.019,-45.236,-118.38,-587.69,0.0000,-1061.9,-1536.7,-748.29,-1211.2
1222.000000000,93.616,2056.5,2119.2,1759.0,311.07,3768.5,969.18,3.1926,6112.1,2716.8,3361.8,2043.7,0.0000,-6579.0,-6874.3,-1318.7,-2122.1,-2064.9,-15712.,-108.93,-19361.,-6176.0,-4077.0,-2417.0,67.544,2406.2,2194.1,1839.4,341.53,4090.3,1686.6,0.0000,7284.3,4449.7,4252.8,3658.0,0.0000,-373.65,-114.39,-97.679,-45.029,-118.08,-587.69,0.0000,-1061.9,-1536.6,-748.28,-1211.1
1223.000000000,93.230,2047.9,2110.3,1755.7,309.74,3765.2,969.18,3.1994,6110.9,2716.7,3362.0,2043.8,0.0000,-6576.6,-6873.0,-1318.5,-2121.3,-2065.0,-15711.,-108.89,-19360.,-6175.6,-4076.5,-2416.2,67.223,2394.8,2183.6,1833.5,339.95,4078.5,1686.6,0.0000,7277.2,4449.7,4252.8,3658.0,0.0000,-371.85,-113.82,-97.311,-44.815,-117.73,-587.69,0.0000,-1061.8,-1536.6,-748.26,-1211.0
1224.000000000,92.734,2039.7,2101.1,1752.0,308.41,3760.5,969.18,3.2105,6110.7,2716.8,3362.2,2043.9,0.0000,-6573.9,-6871.5,-1318.3,-2120.5,-2065.0,-15709.,-108.84,-19359.,-6175.2,-4075.9,-2415.5,66.898,2383.2,2173.1,1827.1,338.35,4065.5,1686.6,0.0000,7269.4,4449.7,4252.8,3658.0,0.0000,-370.02,-113.25,-96.924,-44.598,-117.35,-587.69,0.0000,-1061.7,-1536.5,-748.25,-1210.9
1225.000000000,92.414,2030.9,2092.8,1747.9,307.26,3754.0,969.15,3.2108,6110.7,2716.9,3362.1,2043.9,0.0000,-6570.8,-6869.8,-1318.0,-2119.7,-2064.9,-15708.,-108.80,-19358.,-6174.7,-4075.4,-2414.8,66.660,2374.7,2165.4,1822.6,337.19,4056.6,1686.6,0.0000,7264.0,4449.7,4252.8,3658.0,0.0000,-368.67,-112.82,-96.650,-44.440,-117.08,-587.69,0.0000,-1061.7,-1536.4,-748.23,-1210.7
1226.000000000,92.135,2022.7,2086.0,1743.3,306.12,3748.7,969.15,3.2110,6109.2,2717.1,3362.3,2043.9,0.0000,-6567.5,-6868.0,-1317.6,-2118.9,-2064.7,-15706.,-108.76,-19357.,-6174.3,-4074.9,-2414.1,66.328,2362.9,2154.6,1815.3,335.54,4041.4,1686.6,0.0000,7254.8,4449.7,4252.8,3658.0,0.0000,-366.80,-112.23,-96.230,-44.219,-116.62,-587.69,0.0000,-1061.6,-1536.3,-748.22,-1210.6
1227.000000000,91.990,2014.4,2080.5,1738.3,304.74,3741.8,969.15,3.2113,6107.4,2717.2,3362.4,2044.0,0.0000,-6564.1,-6866.1,-1317.1,-2118.1,-2064.5,-15705.,-108.72,-19356.,-6173.9,-4074.4,-2413.3,65.990,2350.9,2143.6,1807.5,333.85,4025.0,1686.6,0.0000,7244.9,4449.7,4252.8,3658.0,0.0000,-364.88,-111.63,-95.789,-43.993,-116.13,-587.69,0.0000,-1061.5,-1536.2,-748.21,-1210.5
1228.000000000,91.687,2005.4,2071.1,1732.8,303.40,3732.6,969.15,3.2116,6103.1,2717.3,3362.4,2044.0,0.0000,-6560.4,-6864.0,-1316.5,-2117.3,-2064.3,-15703.,-108.67,-19355.,-6173.5,-4073.9,-2412.6,65.659,2339.1,2132.8,1799.6,332.20,4008.0,1686.6,0.0000,7234.7,4449.7,4252.8,3658.0,0.0000,-363.01,-111.03,-95.347,-43.773,-115.62,-587.69,0.0000,-1061.4,-1536.2,-748.19,-1210.4
1229.000000000,91.367,1996.1,2061.5,1728.3,301.90,3722.5,969.16,3.2118,6097.9,2717.6,3362.2,2044.2,0.0000,-6556.5,-6861.7,-1315.8,-2116.4,-2064.0,-15702.,-108.63,-19354.,-6173.0,-4073.3,-2411.9,65.357,2328.3,2123.0,1791.8,330.68,3991.3,1686.6,0.0000,7224.6,4449.7,4252.8,3658.0,0.0000,-361.28,-110.48,-94.926,-43.571,-115.11,-587.69,0.0000,-1061.4,-1536.1,-748.18,-1210.3
1230.000000000,91.047,1986.9,2053.9,1722.5,300.50,3711.4,969.16,3.2121,6092.0,2717.8,3362.1,2044.4,0.0000,-6552.4,-6859.4,-1315.0,-2115.5,-2063.5,-15700.,-108.59,-19353.,-6172.6,-4072.8,-2411.2,65.037,2316.9,2112.6,1783.4,329.06,3973.0,1686.6,0.0000,7213.5,4449.7,4252.8,3658.0,0.0000,-359.46,-109.90,-94.474,-43.358,-114.56,-587.69,0.0000,-1061.3,-1536.0,-748.16,-1210.2
1231.000000000,90.659,1978.9,2047.3,1716.1,299.31,3700.7,969.16,3.2123,6085.7,2717.8,3362.1,2044.5,0.0000,-6548.1,-6857.0,-1314.2,-2114.5,-2062.9,-15699.,-108.55,-19351.,-6172.2,-4072.3,-2410.4,64.987,2336.0,2111.0,1779.4,328.76,3962.0,1686.6,0.0000,7206.8,4449.7,4252.8,3658.0,0.0000,-359.16,-109.78,-94.295,-43.325,-114.21,-587.69,0.0000,-1061.2,-1535.9,-748.15,-1210.0
1232.000000000,90.268,1973.3,2041.0,1709.7,298.54,3689.7,969.16,3.2122,6079.0,2717.8,3362.1,2044.6,0.0000,-6543.9,-6854.7,-1313.3,-2113.6,-2062.2,-15697.,-108.50,-19350.,-6171.8,-4071.8,-2409.7,64.805,2308.7,2105.1,1773.1,327.83,3949.0,1686.6,0.0000,7198.9,4449.7,4252.8,3658.0,0.0000,-358.07,-109.43,-94.003,-43.204,-113.80,-587.69,0.0000,-1061.1,-1535.8,-748.14,-1209.9
1233.000000000,90.060,1967.4,2034.3,1703.7,297.55,3679.4,969.16,3.2208,6072.1,2717.9,3361.9,2044.6,0.0000,-6539.6,-6852.4,-1312.3,-2112.7,-2061.4,-15696.,-108.46,-19349.,-6171.4,-4071.3,-2409.0,64.512,2298.2,2095.6,1764.4,326.33,3929.6,1686.6,0.0000,7187.2,4449.7,4252.8,3658.0,0.0000,-356.39,-108.90,-93.554,-43.008,-113.20,-587.69,0.0000,-1061.0,-1535.8,-748.12,-1209.8
1234.000000000,89.819,1962.4,2028.8,1697.8,296.97,3667.9,969.16,3.2255,6066.0,2718.0,3362.0,2044.7,0.0000,-6535.3,-6850.1,-1311.4,-2111.8,-2060.6,-15694.,-108.42,-19348.,-6171.0,-4070.8,-2408.3,89.887,2315.6,2136.9,1764.5,335.41,3926.7,1686.6,0.0000,7185.4,4449.7,4252.8,3658.0,0.0000,-357.85,-110.02,-93.697,-43.239,-113.09,-587.69,0.0000,-1061.0,-1535.7,-748.11,-1209.7
1235.000000000,89.782,1966.3,2031.3,1692.8,297.86,3660.0,969.16,2.5040,6059.1,2718.1,3362.0,2044.8,0.0000,-6531.7,-6848.2,-1310.5,-2111.0,-2059.7,-15692.,-108.38,-19347.,-6170.6,-4070.2,-2407.6,183.09,2400.8,2298.8,1784.1,357.33,3960.2,1686.6,43.931,7207.9,4459.9,4264.4,3672.4,0.0000,-363.15,-114.39,-94.681,-43.981,-113.87,-587.69,-2.0058,-1061.2,-1535.6,-748.15,-1209.9
1236.000000000,90.182,1979.3,2042.5,1691.5,299.77,3657.1,969.16,2.2708,6054.2,2718.2,3362.1,2044.9,0.0000,-6529.3,-6847.1,-1309.7,-2110.3,-2059.0,-15691.,-108.34,-19346.,-6170.2,-4069.7,-2406.8,66.199,2362.8,2150.4,1778.1,334.31,3946.3,1686.6,0.0000,7197.0,4449.7,4252.8,3658.0,0.0000,-365.55,-111.66,-94.890,-44.133,-113.59,-587.69,0.0000,-1061.0,-1535.5,-748.08,-1209.5
1237.000000000,90.649,1989.0,2051.9,1692.1,301.17,3653.1,969.17,2.2711,6049.6,2718.3,3362.1,2045.1,0.0000,-6527.5,-6846.4,-1309.0,-2109.7,-2058.3,-15689.,-108.30,-19345.,-6169.8,-4069.2,-2406.1,66.141,2356.3,2148.5,1770.1,333.91,3926.0,1686.6,0.0000,7184.7,4449.7,4252.8,3658.0,0.0000,-365.19,-111.54,-94.586,-44.094,-112.97,-587.69,0.0000,-1060.9,-1535.5,-748.07,-1209.4
1238.000000000,90.976,1990.9,2054.5,1691.1,301.95,3645.4,969.12,2.2713,6044.3,2718.2,3362.1,2045.2,0.0000,-6525.8,-6845.6,-1308.3,-2109.1,-2057.5,-15688.,-108.26,-19343.,-6169.3,-4068.7,-2405.4,65.957,2349.7,2142.5,1760.9,332.90,3904.2,1686.6,0.0000,7171.5,4449.7,4252.8,3658.0,0.0000,-364.13,-111.21,-94.176,-43.971,-112.30,-587.69,0.0000,-1060.8,-1535.4,-748.05,-1209.2
1239.000000000,91.110,1988.3,2052.7,1687.3,301.79,3636.0,969.12,2.2716,6039.2,2718.3,3362.2,2045.3,0.0000,-6523.9,-6844.6,-1307.5,-2108.4,-2056.5,-15686.,-108.22,-19342.,-6168.9,-4068.2,-2404.7,65.720,2341.3,2134.8,1751.3,331.65,3882.0,1686.6,0.0000,7158.0,4449.7,4252.8,3658.0,0.0000,-362.79,-110.79,-93.726,-43.814,-111.61,-587.69,0.0000,-1060.7,-1535.3,-748.04,-1209.1
1240.000000000,91.124,1983.5,2048.1,1681.5,300.87,3622.8,969.12,2.2718,6034.5,2718.5,3362.2,2045.4,0.0000,-6521.6,-6843.5,-1306.6,-2107.6,-2055.4,-15685.,-108.18,-19341.,-6168.5,-4067.7,-2404.0,65.452,2331.7,2126.1,1741.4,330.25,3859.3,1686.6,0.0000,7144.3,4449.7,4252.8,3658.0,0.0000,-361.27,-110.32,-93.249,-43.635,-110.91,-587.69,0.0000,-1060.6,-1535.2,-748.03,-1209.0
1241.000000000,90.840,1977.4,2042.5,1674.2,299.75,3609.9,969.12,1.9651,6031.2,2718.6,3362.3,2045.5,0.0000,-6518.8,-6842.1,-1305.5,-2106.8,-2054.1,-15683.,-108.14,-19339.,-6168.1,-4067.2,-2403.3,65.167,2321.5,2116.8,1731.3,328.77,3836.2,1686.6,0.0000,7130.3,4449.7,4252.8,3658.0,0.0000,-359.65,-109.81,-92.756,-43.444,-110.20,-587.69,0.0000,-1060.5,-1535.1,-748.01,-1208.9
1242.000000000,90.640,1970.6,2036.4,1665.7,298.51,3598.4,969.13,1.9901,6026.8,2718.7,3362.3,2045.6,0.0000,-6515.8,-6840.6,-1304.3,-2106.0,-2052.6,-15682.,-108.09,-19338.,-6167.7,-4066.7,-2402.6,64.870,2311.0,2107.2,1721.1,327.23,3813.0,1686.6,0.0000,7116.2,4449.7,4252.8,3658.0,0.0000,-357.97,-109.29,-92.253,-43.247,-109.47,-587.69,0.0000,-1060.4,-1535.1,-748.00,-1208.8
1243.000000000,90.594,1963.7,2030.4,1657.3,297.21,3585.1,969.13,2.3446,6019.9,2718.8,3362.3,2045.7,0.0000,-6512.5,-6838.8,-1302.9,-2105.2,-2051.1,-15680.,-108.05,-19337.,-6167.3,-4066.2,-2401.8,64.575,2300.5,2097.6,1710.8,325.70,3789.5,1686.6,0.0000,7102.0,4449.7,4252.8,3658.0,0.0000,-356.29,-108.76,-91.749,-43.050,-108.74,-587.69,0.0000,-1060.3,-1535.0,-747.98,-1208.7
1244.000000000,90.349,1956.3,2022.5,1649.8,295.89,3568.2,969.13,2.3448,6010.7,2718.8,3362.3,2045.8,0.0000,-6508.9,-6837.0,-1301.5,-2104.3,-2049.4,-15678.,-108.01,-19335.,-6166.9,-4065.7,-2401.1,64.277,2289.8,2088.0,1700.5,324.16,3766.3,1686.6,0.0000,7088.0,4449.7,4252.8,3658.0,0.0000,-354.60,-108.23,-91.246,-42.852,-108.01,-587.69,0.0000,-1060.2,-1534.9,-747.97,-1208.6
1245.000000000,90.051,1948.5,2014.0,1641.6,294.55,3549.3,969.13,2.3589,6000.0,2718.8,3362.2,2045.9,0.0000,-6504.9,-6835.0,-1300.0,-2103.4,-2047.6,-15677.,-107.97,-19334.,-6166.5,-4065.2,-2400.4,63.982,2279.3,2078.4,1690.4,322.63,3743.2,1686.6,0.0000,7074.0,4449.7,4252.8,3658.0,0.0000,-352.91,-107.70,-90.746,-42.655,-107.29,-587.69,0.0000,-1060.0,-1534.8,-747.96,-1208.5
1246.000000000,90.021,1941.4,2005.9,1632.7,293.25,3530.0,969.13,2.3599,5988.5,2718.9,3362.2,2046.0,0.0000,-6500.6,-6832.9,-1298.4,-2102.5,-2045.7,-15675.,-107.93,-19332.,-6166.1,-4064.7,-2399.7,63.733,2270.4,2070.3,1680.9,321.32,3721.5,1686.6,0.0000,7060.9,4449.7,4252.8,3658.0,0.0000,-351.48,-107.24,-90.294,-42.489,-106.60,-587.69,0.0000,-1059.9,-1534.7,-747.94,-1208.3
1247.000000000,89.750,1934.3,1998.1,1623.7,292.00,3511.3,969.13,2.3601,5977.2,2718.9,3362.2,2046.1,0.0000,-6496.1,-6830.7,-1296.8,-2101.6,-2043.8,-15674.,-107.89,-19331.,-6165.7,-4064.2,-2399.0,63.439,2260.0,2060.7,1670.7,319.80,3698.3,1686.6,0.0000,7046.8,4449.7,4252.8,3658.0,0.0000,-349.80,-106.71,-89.795,-42.293,-105.86,-587.69,0.0000,-1059.8,-1534.7,-747.93,-1208.2
1248.000000000,89.515,1927.4,1990.4,1615.3,290.76,3492.6,969.13,2.3604,5966.0,2719.0,3362.2,2046.2,0.0000,-6491.3,-6828.5,-1295.1,-2100.6,-2041.8,-15672.,-107.84,-19329.,-6165.3,-4063.6,-2398.3,63.232,2252.6,2054.0,1661.8,318.70,3677.4,1686.6,0.0000,7034.2,4449.7,4252.8,3658.0,0.0000,-348.59,-106.32,-89.382,-42.155,-105.19,-587.69,0.0000,-1059.7,-1534.6,-747.92,-1208.1
1249.000000000,89.117,1929.5,1990.6,1607.8,291.01,3477.5,969.13,2.3607,5954.8,2719.1,3362.2,2046.3,0.0000,-6487.1,-6826.6,-1293.5,-2099.8,-2039.8,-15671.,-107.81,-19328.,-6164.9,-4063.1,-2397.6,132.07,2370.9,2217.8,1702.0,337.65,3757.8,1686.6,89.847,7085.0,4456.8,4260.4,3666.4,0.0000,-357.09,-111.30,-91.366,-43.246,-107.31,-587.69,-4.1023,-1060.0,-1534.5,-747.94,-1208.2
1250.000000000,89.649,1947.2,2004.9,1606.6,294.00,3473.5,969.13,2.3610,5946.6,2719.1,3362.2,2046.5,0.0000,-6484.5,-6825.7,-1292.2,-2099.1,-2038.0,-15669.,-107.77,-19326.,-6164.5,-4062.6,-2396.8,96.350,2452.4,2379.6,1715.6,366.32,3784.3,1686.6,54.182,7098.7,4482.7,4305.0,3722.7,0.0000,-360.62,-115.36,-91.882,-43.825,-107.56,-587.69,-2.4739,-1060.1,-1534.4,-748.15,-1209.1
1251.000000000,90.024,1963.7,2020.8,1611.0,296.08,3473.9,969.13,2.3613,5941.1,2719.1,3362.3,2046.6,0.0000,-6483.1,-6825.5,-1291.2,-2098.5,-2036.6,-15667.,-107.73,-19324.,-6164.1,-4062.1,-2396.1,65.794,2343.9,2137.2,1700.8,333.11,3759.8,1686.6,0.0000,7084.9,4474.7,4296.5,3707.1,0.0000,-362.58,-110.57,-91.956,-43.875,-107.03,-587.69,0.0000,-1060.0,-1534.4,-748.09,-1208.7
1252.000000000,90.554,1973.8,2030.4,1614.0,298.37,3469.3,969.14,2.3616,5935.0,2719.1,3362.3,2046.7,0.0000,-6482.2,-6825.6,-1290.2,-2098.0,-2035.3,-15666.,-107.69,-19323.,-6163.7,-4061.6,-2395.4,65.733,2341.7,2135.3,1691.7,331.17,3731.1,1686.6,0.0000,7066.7,4459.8,4268.9,3675.2,0.0000,-362.22,-110.46,-91.667,-43.825,-106.39,-587.69,0.0000,-1059.8,-1534.3,-747.94,-1208.0
1253.000000000,90.967,1976.3,2033.9,1614.6,299.02,3460.3,969.14,2.3619,5927.6,2719.1,3362.3,2046.8,0.0000,-6481.3,-6825.5,-1289.1,-2097.4,-2033.7,-15664.,-107.65,-19321.,-6163.3,-4061.1,-2394.7,65.585,2336.4,2130.4,1683.0,329.91,3707.1,1686.6,0.0000,7051.9,4452.1,4256.8,3662.2,0.0000,-361.37,-110.20,-91.313,-43.723,-105.75,-587.69,0.0000,-1059.7,-1534.2,-747.87,-1207.6
1254.000000000,91.209,1975.2,2033.1,1612.0,298.89,3448.1,969.14,1.8983,5921.5,2719.0,3362.3,2046.8,0.0000,-6480.0,-6825.1,-1288.2,-2096.8,-2032.0,-15662.,-107.61,-19319.,-6162.9,-4060.6,-2394.0,65.382,2329.2,2123.9,1674.3,328.78,3685.8,1686.6,0.0000,7038.9,4450.1,4253.4,3658.5,0.0000,-360.23,-109.85,-90.913,-43.588,-105.10,-587.69,0.0000,-1059.5,-1534.1,-747.84,-1207.5
1255.000000000,91.162,1971.6,2029.7,1607.3,298.15,3434.9,969.14,2.1555,5918.3,2719.2,3362.4,2046.9,0.0000,-6478.4,-6824.6,-1287.1,-2096.1,-2030.1,-15661.,-107.57,-19318.,-6162.5,-4060.1,-2393.3,65.148,2320.9,2116.2,1665.3,327.55,3664.9,1686.6,0.0000,7026.2,4449.7,4252.8,3658.0,0.0000,-358.91,-109.44,-90.485,-43.432,-104.44,-587.69,0.0000,-1059.4,-1534.1,-747.82,-1207.3
1256.000000000,90.812,1966.5,2025.9,1600.5,297.17,3426.5,969.14,2.4315,5920.2,2719.3,3362.5,2047.0,0.0000,-6476.4,-6823.8,-1285.8,-2095.4,-2028.0,-15659.,-107.53,-19316.,-6162.1,-4059.6,-2392.6,64.889,2311.7,2107.8,1656.0,326.20,3643.6,1686.6,0.0000,7013.3,4449.7,4252.8,3658.0,0.0000,-357.45,-108.99,-90.034,-43.260,-103.76,-587.69,0.0000,-1059.3,-1534.0,-747.81,-1207.2
1257.000000000,90.581,1961.1,2021.5,1592.7,296.05,3419.6,969.14,2.4318,5917.7,2719.4,3362.6,2047.1,0.0000,-6474.1,-6822.7,-1284.4,-2094.7,-2025.9,-15658.,-107.49,-19314.,-6161.7,-4059.1,-2391.9,64.618,2302.0,2099.0,1646.5,324.80,3622.1,1686.6,0.0000,7000.2,4449.7,4252.8,3658.0,0.0000,-355.92,-108.52,-89.571,-43.079,-103.08,-587.69,0.0000,-1059.2,-1533.9,-747.79,-1207.1
1258.000000000,90.327,1954.9,2016.5,1586.5,294.85,3407.3,969.14,2.4321,5911.8,2719.4,3362.6,2047.1,0.0000,-6471.6,-6821.5,-1282.8,-2093.9,-2023.7,-15656.,-107.45,-19313.,-6161.3,-4058.6,-2391.2,64.338,2292.0,2089.9,1636.9,323.35,3600.3,1686.6,0.0000,6987.0,4449.7,4252.8,3658.0,0.0000,-354.34,-108.02,-89.098,-42.892,-102.38,-587.69,0.0000,-1059.1,-1533.8,-747.78,-1207.0
1259.000000000,90.056,1948.0,2010.3,1580.1,293.62,3390.9,969.14,2.4324,5902.9,2719.3,3362.6,2047.2,0.0000,-6468.7,-6820.2,-1281.2,-2093.0,-2021.4,-15654.,-107.40,-19311.,-6160.9,-4058.1,-2390.4,64.056,2282.0,2080.8,1627.3,321.89,3578.5,1686.6,0.0000,6973.8,4449.7,4252.8,3658.0,0.0000,-352.74,-107.52,-88.623,-42.704,-101.68,-587.69,0.0000,-1059.0,-1533.8,-747.76,-1206.9
1260.000000000,89.778,1941.6,2002.9,1572.5,292.39,3374.3,969.14,2.4326,5892.2,2719.3,3362.7,2047.2,0.0000,-6465.4,-6818.7,-1279.6,-2092.2,-2019.0,-15653.,-107.36,-19309.,-6160.4,-4057.6,-2389.7,63.815,2273.4,2072.9,1617.9,320.62,3556.8,1686.6,0.0000,6960.7,4449.7,4252.8,3658.0,0.0000,-351.37,-107.09,-88.178,-42.543,-100.99,-587.69,0.0000,-1058.9,-1533.7,-747.75,-1206.8
1261.000000000,89.516,1935.2,1995.7,1564.1,291.12,3356.9,969.14,2.5049,5880.9,2719.3,3362.7,2047.3,0.0000,-6461.9,-6817.1,-1277.9,-2091.4,-2016.5,-15651.,-107.32,-19307.,-6160.0,-4057.1,-2389.0,63.515,2262.7,2063.2,1607.9,319.07,3534.2,1686.6,0.0000,6947.0,4449.7,4252.8,3658.0,0.0000,-349.66,-106.56,-87.680,-42.343,-100.26,-587.69,0.0000,-1058.8,-1533.6,-747.74,-1206.7
1262.000000000,89.229,1927.6,1988.4,1555.7,289.81,3339.5,969.15,3.1204,5870.4,2719.2,3362.7,2047.4,0.0000,-6458.0,-6815.3,-1276.1,-2090.5,-2014.0,-15649.,-107.28,-19305.,-6159.6,-4056.6,-2388.3,63.216,2252.1,2053.5,1597.9,317.53,3511.5,1686.6,0.0000,6933.3,4449.7,4252.8,3658.0,0.0000,-347.97,-106.03,-87.185,-42.144,-99.534,-587.69,0.0000,-1058.6,-1533.5,-747.72,-1206.6
1263.000000000,88.939,1919.8,1981.0,1547.1,288.51,3323.0,969.15,3.1207,5859.6,2719.2,3362.7,2047.5,0.0000,-6453.9,-6813.5,-1274.3,-2089.6,-2011.4,-15648.,-107.24,-19304.,-6159.2,-4056.1,-2387.6,62.918,2241.4,2043.8,1587.8,315.99,3488.8,1686.6,0.0000,6919.5,4449.7,4252.8,3658.0,0.0000,-346.27,-105.49,-86.688,-41.945,-98.803,-587.69,0.0000,-1058.5,-1533.5,-747.71,-1206.5
1264.000000000,88.649,1911.8,1973.9,1538.6,287.18,3304.9,969.15,3.1210,5847.9,2719.4,3362.6,2047.6,0.0000,-6449.6,-6811.5,-1272.4,-2088.7,-2008.7,-15646.,-107.20,-19302.,-6158.8,-4055.6,-2386.9,62.623,2230.9,2034.2,1577.9,314.46,3466.3,1686.6,0.0000,6905.9,4449.7,4252.8,3658.0,0.0000,-344.59,-104.96,-86.195,-41.749,-98.075,-587.69,0.0000,-1058.4,-1533.4,-747.70,-1206.3
1265.000000000,88.350,1903.8,1965.7,1529.6,285.85,3285.7,969.15,3.1213,5836.5,2719.5,3362.7,2047.8,0.0000,-6445.1,-6809.4,-1270.5,-2087.8,-2005.9,-15644.,-107.16,-19300.,-6158.4,-4055.1,-2386.2,62.329,2220.4,2024.7,1567.9,312.94,3443.6,1686.6,0.0000,6892.2,4449.7,4252.8,3658.0,0.0000,-342.90,-104.43,-85.702,-41.552,-97.343,-587.69,0.0000,-1058.3,-1533.3,-747.68,-1206.2
1266.000000000,88.052,1895.7,1957.4,1520.4,284.51,3265.9,969.15,3.1307,5825.4,2719.5,3362.7,2047.9,0.0000,-6440.4,-6807.2,-1268.6,-2086.8,-2003.1,-15643.,-107.12,-19298.,-6157.9,-4054.6,-2385.5,62.033,2209.9,2015.1,1557.8,311.41,3420.9,1686.6,0.0000,6878.4,4449.7,4252.8,3658.0,0.0000,-341.21,-103.90,-85.206,-41.356,-96.607,-587.69,0.0000,-1058.2,-1533.2,-747.67,-1206.1
1267.000000000,87.754,1888.6,1949.9,1511.4,283.38,3248.5,969.15,3.2875,5814.1,2719.6,3362.7,2048.0,0.0000,-6435.5,-6805.0,-1266.6,-2085.9,-2000.3,-15641.,-107.08,-19296.,-6157.5,-4054.1,-2384.8,65.287,2209.3,2018.6,1558.1,318.72,3431.0,1686.6,0.0000,6876.7,4449.7,4264.6,3671.1,0.0000,-341.05,-103.92,-85.157,-41.389,-96.506,-587.69,0.0000,-1058.1,-1533.2,-747.72,-1206.3
1268.000000000,87.592,1883.4,1943.9,1503.6,282.61,3231.6,969.15,3.7966,5803.0,2719.7,3362.7,2048.1,0.0000,-6430.6,-6802.7,-1264.7,-2084.9,-1997.4,-15639.,-107.04,-19294.,-6157.1,-4053.6,-2384.1,61.752,2199.9,2005.9,1547.4,309.95,3397.0,1686.6,0.0000,6864.0,4449.7,4252.8,3658.0,0.0000,-339.53,-103.35,-84.706,-41.168,-95.760,-587.69,0.0000,-1058.0,-1533.1,-747.64,-1205.9
1269.000000000,87.360,1877.1,1937.2,1496.9,281.52,3215.2,969.15,3.2720,5792.1,2719.9,3362.7,2048.2,0.0000,-6425.6,-6800.5,-1262.8,-2084.0,-1994.6,-15637.,-107.00,-19292.,-6156.7,-4053.1,-2383.3,61.483,2190.3,1997.2,1537.9,308.55,3375.2,1686.6,0.0000,6850.7,4449.7,4252.8,3658.0,0.0000,-337.99,-102.86,-84.240,-40.989,-95.048,-587.69,0.0000,-1057.9,-1533.0,-747.63,-1205.8
1270.000000000,87.114,1869.8,1929.4,1489.4,280.52,3198.2,969.15,3.1431,5781.6,2720.0,3362.7,2048.3,0.0000,-6420.5,-6798.2,-1260.8,-2083.0,-1991.7,-15636.,-106.96,-19290.,-6156.3,-4052.6,-2382.6,61.212,2180.6,1988.4,1528.1,307.13,3353.0,1686.6,0.0000,6837.3,4449.7,4252.8,3658.0,0.0000,-336.42,-102.36,-83.768,-40.808,-94.327,-587.69,0.0000,-1057.8,-1532.9,-747.61,-1205.7
1271.000000000,86.896,1862.3,1921.3,1481.9,279.36,3179.7,969.15,3.1441,5771.5,2720.1,3362.9,2048.4,0.0000,-6415.2,-6795.8,-1258.9,-2082.0,-1988.7,-15634.,-106.91,-19288.,-6155.9,-4052.1,-2381.9,60.942,2171.0,1979.6,1518.5,305.73,3330.9,1686.6,0.0000,6823.9,4449.7,4252.8,3658.0,0.0000,-334.86,-101.87,-83.298,-40.628,-93.607,-587.69,0.0000,-1057.7,-1532.9,-747.60,-1205.6
1272.000000000,86.693,1854.5,1913.8,1473.6,278.14,3161.2,969.15,3.1492,5760.7,2720.2,3363.0,2048.4,0.0000,-6409.7,-6793.3,-1257.0,-2081.0,-1985.6,-15632.,-106.87,-19286.,-6155.5,-4051.5,-2381.2,60.677,2161.6,1971.0,1508.9,304.35,3309.0,1686.6,0.0000,6810.6,4449.7,4252.8,3658.0,0.0000,-333.33,-101.38,-82.833,-40.451,-92.890,-587.69,0.0000,-1057.5,-1532.8,-747.59,-1205.5
1273.000000000,86.626,1848.3,1908.1,1465.3,277.20,3143.0,969.13,3.1394,5750.0,2720.3,3363.0,2048.5,0.0000,-6404.2,-6790.8,-1255.0,-2080.0,-1982.5,-15631.,-106.83,-19284.,-6155.1,-4051.0,-2380.5,65.530,2172.7,1983.8,1509.5,311.44,3311.9,1686.6,11.028,6809.1,4451.4,4259.2,3664.7,0.0000,-333.94,-101.73,-82.842,-40.573,-92.682,-587.69,-0.50352,-1057.5,-1532.7,-747.61,-1205.5
1274.000000000,86.546,1885.7,1942.0,1459.3,283.51,3133.3,969.11,3.1180,5741.4,2720.4,3363.0,2048.7,0.0000,-6401.9,-6790.2,-1253.7,-2079.4,-1979.5,-15629.,-106.80,-19282.,-6154.7,-4050.5,-2379.8,297.11,2666.0,2604.1,1613.1,368.04,3484.0,1687.5,164.19,6907.2,4460.4,4278.0,3685.1,0.0000,-381.23,-123.35,-90.517,-46.376,-97.001,-587.70,-7.4968,-1058.1,-1532.7,-747.69,-1205.7
1275.000000000,90.770,1996.2,2036.3,1464.8,300.99,3143.3,969.11,2.5030,5737.2,2720.5,3363.0,2048.8,0.0000,-6407.5,-6794.2,-1252.8,-2079.7,-1977.0,-15627.,-106.76,-19280.,-6154.3,-4050.0,-2379.1,71.616,2551.3,2326.3,1630.5,647.77,3531.5,1686.8,0.0000,6898.0,4452.9,4287.4,3673.3,0.0000,-393.37,-119.70,-91.819,-49.541,-96.763,-587.69,0.0000,-1058.0,-1532.6,-747.72,-1205.4
1276.000000000,93.151,2072.6,2115.5,1484.3,308.79,3155.0,969.11,2.5001,5734.8,2720.5,3363.0,2048.9,0.0000,-6416.8,-6800.8,-1252.2,-2080.3,-1975.0,-15625.,-106.73,-19278.,-6153.9,-4049.5,-2378.4,71.763,2556.5,2331.1,1610.1,363.12,3456.5,1686.8,0.0000,6880.2,4450.5,4266.4,3663.2,0.0000,-394.25,-120.02,-91.664,-47.881,-95.882,-587.69,0.0000,-1057.8,-1532.5,-747.60,-1205.1
1277.000000000,94.895,2102.1,2149.2,1497.8,317.76,3156.6,969.09,2.5004,5730.9,2720.6,3363.0,2049.1,0.0000,-6426.3,-6806.7,-1251.7,-2080.8,-1973.1,-15624.,-106.69,-19276.,-6153.5,-4049.0,-2377.7,71.622,2551.5,2326.5,1595.0,357.02,3412.4,1686.8,0.0000,6865.3,4449.9,4256.9,3659.1,0.0000,-393.55,-119.86,-91.294,-47.754,-95.101,-587.69,0.0000,-1057.6,-1532.4,-747.54,-1204.9
1278.000000000,96.842,2111.7,2163.8,1504.3,320.68,3150.3,969.09,2.5008,5724.1,2720.8,3362.9,2049.2,0.0000,-6435.2,-6811.6,-1251.0,-2081.1,-1970.8,-15622.,-106.65,-19274.,-6153.0,-4048.5,-2377.0,71.389,2543.2,2319.0,1583.4,354.78,3382.3,1686.8,0.0000,6852.0,4449.7,4253.4,3658.1,0.0000,-392.36,-119.54,-90.866,-47.592,-94.393,-587.69,0.0000,-1057.5,-1532.4,-747.51,-1204.8
1279.000000000,96.970,2115.0,2170.3,1502.0,320.01,3140.3,969.09,2.5011,5719.9,2720.8,3363.0,2049.3,0.0000,-6442.6,-6815.5,-1250.5,-2081.1,-1968.3,-15620.,-106.61,-19272.,-6152.6,-4048.0,-2376.3,71.098,2532.8,2309.5,1573.6,353.29,3359.5,1686.8,0.0000,6839.2,4449.7,4252.8,3658.0,0.0000,-390.84,-119.12,-90.398,-47.399,-93.714,-587.69,0.0000,-1057.4,-1532.3,-747.49,-1204.7
1280.000000000,96.756,2114.2,2169.2,1501.0,318.83,3126.8,969.09,2.5014,5716.8,2720.8,3363.0,2049.5,0.0000,-6448.8,-6818.8,-1249.8,-2081.1,-1965.6,-15618.,-106.57,-19270.,-6152.2,-4047.5,-2375.6,70.775,2521.3,2299.0,1564.0,351.64,3338.3,1686.8,0.0000,6826.4,4449.7,4252.8,3658.0,0.0000,-389.15,-118.64,-89.907,-47.183,-93.038,-587.69,0.0000,-1057.3,-1532.2,-747.48,-1204.6
1281.000000000,96.406,2109.7,2171.7,1493.7,317.41,3120.4,969.10,2.1212,5723.3,2720.8,3363.0,2049.6,0.0000,-6454.2,-6821.4,-1248.8,-2080.9,-1962.8,-15616.,-106.53,-19268.,-6151.8,-4047.0,-2374.9,70.430,2509.0,2287.8,1554.4,349.90,3317.1,1686.8,0.0000,6813.6,4449.7,4252.8,3658.0,0.0000,-387.33,-118.12,-89.400,-46.953,-92.357,-587.69,0.0000,-1057.2,-1532.2,-747.46,-1204.5
1282.000000000,95.890,2108.6,2173.4,1485.2,315.93,3119.4,969.09,1.8487,5725.1,2720.9,3363.0,2049.7,0.0000,-6459.0,-6823.4,-1247.6,-2080.6,-1959.9,-15615.,-106.49,-19266.,-6151.4,-4046.5,-2374.2,70.073,2496.3,2276.2,1544.7,348.09,3296.0,1686.8,0.0000,6800.8,4449.7,4252.8,3658.0,0.0000,-385.43,-117.56,-88.884,-46.715,-91.675,-587.69,0.0000,-1057.1,-1532.1,-747.45,-1204.4
1283.000000000,95.619,2103.9,2167.3,1480.0,314.38,3113.8,969.05,1.8605,5722.3,2720.8,3363.0,2049.8,0.0000,-6463.1,-6825.1,-1246.4,-2080.2,-1956.9,-15613.,-106.45,-19264.,-6151.0,-4046.0,-2373.5,69.714,2483.5,2264.5,1535.0,346.28,3275.0,1686.7,0.0000,6788.1,4449.7,4252.8,3658.0,0.0000,-383.51,-116.99,-88.369,-46.476,-90.997,-587.69,0.0000,-1057.0,-1532.0,-747.44,-1204.3
1284.000000000,95.102,2095.0,2157.3,1476.5,312.82,3098.5,969.05,1.8608,5714.7,2721.0,3363.0,2049.9,0.0000,-6466.0,-6826.2,-1245.2,-2079.9,-1953.8,-15611.,-106.41,-19262.,-6150.6,-4045.5,-2372.8,69.355,2470.7,2252.9,1525.5,344.47,3254.2,1686.7,0.0000,6775.5,4449.7,4252.8,3658.0,0.0000,-381.58,-116.42,-87.858,-46.237,-90.324,-587.69,0.0000,-1056.8,-1531.9,-747.42,-1204.2
1285.000000000,94.630,2091.9,2148.4,1470.0,311.24,3080.6,969.02,1.2764,5705.1,2721.1,3363.0,2050.0,0.0000,-6467.8,-6827.1,-1243.9,-2079.4,-1950.6,-15609.,-106.37,-19260.,-6150.2,-4045.0,-2372.1,68.998,2458.0,2241.3,1516.0,342.67,3233.6,1686.6,0.0000,6763.1,4449.7,4252.8,3658.0,0.0000,-379.65,-115.84,-87.350,-45.999,-89.655,-587.69,0.0000,-1056.7,-1531.9,-747.41,-1204.1
1286.000000000,94.270,2085.3,2143.2,1461.3,309.67,3062.7,969.00,1.2436,5694.2,2721.0,3363.0,2050.1,0.0000,-6468.8,-6827.8,-1242.6,-2078.9,-1947.4,-15608.,-106.33,-19258.,-6149.8,-4044.4,-2371.4,68.643,2445.4,2229.8,1506.6,340.87,3213.1,1686.6,0.0000,6750.7,4449.7,4252.8,3658.0,0.0000,-377.72,-115.26,-86.844,-45.762,-88.990,-587.69,0.0000,-1056.6,-1531.8,-747.40,-1204.0
1287.000000000,93.912,2075.3,2134.3,1452.5,308.15,3045.7,968.98,1.3214,5683.5,2721.0,3362.9,2050.2,0.0000,-6469.1,-6828.1,-1241.2,-2078.4,-1944.1,-15606.,-106.29,-19256.,-6149.4,-4043.9,-2370.7,68.293,2432.9,2218.4,1497.2,339.11,3192.8,1686.6,0.0000,6738.4,4449.7,4252.8,3658.0,0.0000,-375.81,-114.68,-86.345,-45.528,-88.329,-587.69,0.0000,-1056.5,-1531.7,-747.38,-1203.8
1288.000000000,93.556,2068.5,2126.0,1443.8,306.72,3030.9,968.98,1.9184,5674.2,2721.0,3362.9,2050.3,0.0000,-6469.1,-6828.3,-1239.7,-2077.9,-1940.9,-15604.,-106.25,-19254.,-6149.0,-4043.4,-2370.0,67.943,2420.4,2207.0,1488.0,337.34,3172.6,1686.6,0.0000,6726.2,4449.7,4252.8,3658.0,0.0000,-373.90,-114.10,-85.840,-45.295,-87.671,-587.69,0.0000,-1056.4,-1531.7,-747.37,-1203.7
1289.000000000,93.203,2058.5,2121.7,1435.5,305.21,3016.8,968.98,1.9187,5663.9,2721.1,3362.9,2050.4,0.0000,-6468.9,-6828.2,-1238.2,-2077.3,-1937.6,-15602.,-106.21,-19251.,-6148.6,-4042.9,-2369.3,67.594,2408.0,2195.7,1478.7,335.58,3152.5,1686.6,0.0000,6714.1,4449.7,4252.8,3658.0,0.0000,-371.98,-113.51,-85.335,-45.063,-87.013,-587.69,0.0000,-1056.3,-1531.6,-747.36,-1203.6
1290.000000000,92.812,2050.5,2111.4,1427.8,303.72,2999.3,968.98,1.9190,5652.7,2721.2,3362.9,2050.5,0.0000,-6468.2,-6827.8,-1236.6,-2076.7,-1934.2,-15600.,-106.17,-19249.,-6148.2,-4042.4,-2368.7,67.248,2395.7,2184.5,1469.5,333.84,3132.4,1686.6,0.0000,6701.9,4449.7,4252.8,3658.0,0.0000,-370.07,-112.93,-84.832,-44.832,-86.358,-587.69,0.0000,-1056.2,-1531.5,-747.34,-1203.5
1291.000000000,92.423,2041.5,2101.5,1419.4,302.20,2981.3,968.94,1.9193,5641.9,2721.3,3362.9,2050.6,0.0000,-6467.0,-6827.2,-1235.0,-2076.1,-1930.8,-15599.,-106.13,-19247.,-6147.8,-4041.9,-2368.0,66.903,2383.4,2173.2,1460.3,332.10,3112.4,1686.6,0.0000,6689.9,4449.7,4252.8,3658.0,0.0000,-368.17,-112.34,-84.330,-44.602,-85.704,-587.69,0.0000,-1056.1,-1531.4,-747.33,-1203.4
1292.000000000,92.074,2031.2,2091.3,1410.8,300.68,2963.1,968.90,1.9196,5632.1,2721.4,3362.9,2050.7,0.0000,-6465.2,-6826.3,-1233.3,-2075.4,-1927.4,-15597.,-106.09,-19245.,-6147.4,-4041.4,-2367.3,66.563,2371.3,2162.2,1451.2,330.38,3092.6,1686.6,0.0000,6677.9,4449.7,4252.8,3658.0,0.0000,-366.29,-111.75,-83.834,-44.375,-85.054,-587.69,0.0000,-1055.9,-1531.4,-747.31,-1203.3
1293.000000000,91.681,2021.1,2080.8,1403.5,299.14,2945.8,968.90,1.9200,5621.4,2721.5,3363.0,2050.8,0.0000,-6463.1,-6825.2,-1231.6,-2074.7,-1923.9,-15595.,-106.05,-19243.,-6147.0,-4040.9,-2366.6,66.231,2359.5,2151.4,1442.2,328.70,3073.2,1686.6,0.0000,6666.1,4449.7,4252.8,3658.0,0.0000,-364.44,-111.18,-83.347,-44.154,-84.413,-587.69,0.0000,-1055.8,-1531.3,-747.30,-1203.2
1294.000000000,91.342,2011.1,2070.6,1395.7,297.55,2928.4,968.90,1.9202,5611.0,2721.4,3362.9,2050.9,0.0000,-6460.5,-6823.9,-1229.8,-2073.9,-1920.4,-15593.,-106.01,-19241.,-6146.6,-4040.4,-2365.9,65.905,2347.8,2140.8,1433.4,327.06,3053.8,1686.6,0.0000,6654.4,4449.7,4252.8,3658.0,0.0000,-362.62,-110.61,-82.867,-43.937,-83.777,-587.69,0.0000,-1055.7,-1531.2,-747.29,-1203.1
1295.000000000,90.921,2003.1,2060.7,1387.7,296.11,2910.8,968.91,1.9206,5600.2,2721.5,3363.0,2051.0,0.0000,-6457.6,-6822.4,-1228.0,-2073.2,-1916.9,-15591.,-105.97,-19238.,-6146.2,-4039.8,-2365.2,65.582,2336.3,2130.4,1424.6,325.42,3034.7,1686.6,0.0000,6642.8,4449.7,4252.8,3658.0,0.0000,-360.81,-110.05,-82.390,-43.722,-83.144,-587.69,0.0000,-1055.6,-1531.2,-747.27,-1203.0
1296.000000000,90.565,1993.7,2051.6,1380.9,294.68,2894.3,968.91,1.9209,5589.8,2721.4,3363.0,2051.2,0.0000,-6454.4,-6820.7,-1226.2,-2072.4,-1913.3,-15589.,-105.93,-19236.,-6145.8,-4039.3,-2364.5,65.263,2325.0,2120.0,1415.9,323.81,3015.6,1686.6,0.0000,6631.3,4449.7,4252.8,3658.0,0.0000,-359.02,-109.48,-81.918,-43.509,-82.515,-587.69,0.0000,-1055.5,-1531.1,-747.26,-1202.9
1297.000000000,90.452,1984.4,2042.9,1372.6,293.22,2877.2,968.91,2.1451,5580.4,2721.4,3363.0,2051.3,0.0000,-6450.9,-6818.8,-1224.3,-2071.5,-1909.6,-15588.,-105.89,-19234.,-6145.4,-4038.8,-2363.8,64.949,2313.8,2109.8,1407.3,322.22,2996.8,1686.6,0.0000,6619.9,4449.7,4252.8,3658.0,0.0000,-357.25,-108.93,-81.451,-43.300,-81.891,-587.69,0.0000,-1055.4,-1531.0,-747.25,-1202.7
1298.000000000,90.132,1975.9,2040.6,1364.4,291.76,2860.0,968.91,2.5810,5571.2,2721.4,3363.1,2051.4,0.0000,-6447.4,-6816.7,-1222.5,-2070.7,-1905.9,-15586.,-105.85,-19232.,-6144.9,-4038.3,-2363.1,64.640,2302.8,2099.7,1398.7,320.65,2978.1,1686.6,0.0000,6608.6,4449.7,4252.8,3658.0,0.0000,-355.50,-108.37,-80.989,-43.093,-81.270,-587.69,0.0000,-1055.3,-1531.0,-747.23,-1202.6
1299.000000000,89.816,1967.6,2031.2,1356.2,290.39,2844.5,968.91,2.5813,5560.5,2721.5,3363.1,2051.5,0.0000,-6443.7,-6814.6,-1220.5,-2069.9,-1902.2,-15584.,-105.81,-19229.,-6144.5,-4037.8,-2362.4,64.330,2291.7,2089.7,1390.2,319.09,2959.3,1686.6,0.0000,6597.3,4449.7,4252.8,3658.0,0.0000,-353.75,-107.82,-80.527,-42.887,-80.650,-587.69,0.0000,-1055.2,-1530.9,-747.22,-1202.5
1300.000000000,89.502,1958.3,2021.5,1348.1,289.03,2828.0,968.91,2.5816,5550.6,2721.7,3363.1,2051.6,0.0000,-6439.8,-6812.3,-1218.6,-2069.0,-1898.5,-15582.,-105.77,-19227.,-6144.1,-4037.3,-2361.7,64.023,2280.8,2079.7,1381.7,317.53,2940.7,1686.6,0.0000,6586.0,4449.7,4252.8,3658.0,0.0000,-352.01,-107.27,-80.069,-42.682,-80.032,-587.69,0.0000,-1055.1,-1530.8,-747.21,-1202.4
1301.000000000,88.976,1949.3,2013.6,1341.8,287.68,2811.3,968.88,2.1045,5539.9,2721.7,3363.1,2051.7,0.0000,-6435.8,-6809.9,-1216.6,-2068.1,-1894.7,-15580.,-105.73,-19225.,-6143.7,-4036.8,-2361.0,63.718,2269.9,2069.8,1373.2,315.99,2922.2,1686.6,0.0000,6574.8,4449.7,4252.8,3658.0,0.0000,-350.28,-106.72,-79.612,-42.479,-79.417,-587.69,0.0000,-1055.0,-1530.7,-747.19,-1202.3
1302.000000000,88.681,1940.3,2007.8,1333.8,286.33,2794.3,968.87,1.9264,5529.3,2721.8,3363.1,2051.8,0.0000,-6431.7,-6807.5,-1214.6,-2067.2,-1890.9,-15578.,-105.69,-19222.,-6143.3,-4036.2,-2360.3,63.418,2259.2,2060.0,1364.9,314.47,2903.9,1686.6,0.0000,6563.7,4449.7,4252.8,3658.0,0.0000,-348.57,-106.18,-79.162,-42.279,-78.807,-587.69,0.0000,-1054.9,-1530.7,-747.18,-1202.2
1303.000000000,88.490,1931.1,1999.1,1325.9,285.01,2778.1,968.87,1.9268,5518.9,2721.8,3363.2,2051.9,0.0000,-6427.3,-6804.9,-1212.6,-2066.3,-1887.1,-15576.,-105.65,-19220.,-6142.9,-4035.7,-2359.6,63.130,2249.0,2050.7,1356.7,313.00,2886.0,1686.6,0.0000,6552.9,4449.7,4252.8,3658.0,0.0000,-346.92,-105.65,-78.725,-42.087,-78.210,-587.69,0.0000,-1054.7,-1530.6,-747.16,-1202.1
1304.000000000,88.192,1922.8,1990.6,1318.1,283.81,2761.8,968.87,1.9271,5508.5,2721.9,3363.2,2051.9,0.0000,-6422.9,-6802.3,-1210.6,-2065.3,-1883.2,-15575.,-105.61,-19218.,-6142.5,-4035.2,-2358.9,62.978,2243.6,2045.8,1354.8,313.62,2887.2,1686.6,3.5285,6551.5,4450.9,4256.9,3660.6,0.0000,-346.02,-105.36,-78.549,-41.994,-78.002,-587.69,-0.16111,-1054.7,-1530.5,-747.17,-1202.0
1305.000000000,87.965,1916.1,1983.1,1311.1,282.82,2747.2,968.87,2.1750,5498.4,2722.0,3363.2,2051.9,0.0000,-6418.3,-6799.7,-1208.6,-2064.4,-1879.2,-15573.,-105.57,-19215.,-6142.1,-4034.7,-2358.2,62.736,2234.9,2037.9,1347.2,311.03,2865.7,1686.6,0.0000,6540.6,4449.7,4252.8,3658.0,0.0000,-344.62,-104.91,-78.175,-41.824,-77.447,-587.69,0.0000,-1054.6,-1530.5,-747.14,-1201.9
1306.000000000,87.719,1908.7,1975.6,1304.9,281.77,2732.7,968.88,2.6195,5488.6,2722.1,3363.2,2052.0,0.0000,-6413.5,-6797.1,-1206.6,-2063.4,-1875.3,-15571.,-105.53,-19213.,-6141.7,-4034.2,-2357.5,62.463,2225.2,2029.0,1339.4,309.65,2848.6,1686.6,0.0000,6530.3,4449.7,4252.8,3658.0,0.0000,-343.05,-104.41,-77.760,-41.642,-76.874,-587.69,0.0000,-1054.5,-1530.4,-747.12,-1201.8
1307.000000000,87.494,1900.7,1967.5,1298.3,280.73,2718.7,968.88,2.4043,5479.3,2722.2,3363.3,2052.2,0.0000,-6408.6,-6794.5,-1204.5,-2062.5,-1871.4,-15569.,-105.50,-19211.,-6141.3,-4033.7,-2356.9,62.198,2215.8,2020.4,1331.7,308.30,2831.6,1686.6,0.0000,6520.0,4449.7,4252.8,3658.0,0.0000,-341.53,-103.92,-77.350,-41.466,-76.301,-587.69,0.0000,-1054.4,-1530.3,-747.11,-1201.6
1308.000000000,87.303,1892.9,1959.3,1291.8,279.57,2703.3,968.88,2.0003,5470.5,2722.3,3363.3,2052.3,0.0000,-6403.5,-6791.8,-1202.5,-2061.5,-1867.5,-15567.,-105.46,-19208.,-6140.9,-4033.2,-2356.2,61.926,2206.1,2011.6,1323.9,306.92,2814.4,1686.6,0.0000,6509.6,4449.7,4252.8,3658.0,0.0000,-339.96,-103.42,-76.934,-41.284,-75.725,-587.69,0.0000,-1054.3,-1530.3,-747.10,-1201.5
1309.000000000,87.036,1884.9,1951.0,1284.9,278.37,2687.9,968.88,2.0006,5460.7,2722.3,3363.3,2052.4,0.0000,-6398.3,-6789.1,-1200.4,-2060.5,-1863.5,-15565.,-105.42,-19206.,-6140.5,-4032.6,-2355.5,61.649,2196.2,2002.6,1316.0,305.51,2797.0,1686.6,0.0000,6499.1,4449.7,4252.8,3658.0,0.0000,-338.36,-102.91,-76.511,-41.099,-75.143,-587.69,0.0000,-1054.2,-1530.2,-747.08,-1201.4
1310.000000000,86.647,1876.7,1942.5,1277.9,277.09,2673.2,968.88,1.9651,5451.7,2722.4,3363.4,2052.5,0.0000,-6392.9,-6786.3,-1198.3,-2059.5,-1859.4,-15563.,-105.38,-19204.,-6140.1,-4032.1,-2354.8,61.376,2186.5,1993.7,1308.2,304.12,2779.7,1686.6,0.0000,6488.7,4449.7,4252.8,3658.0,0.0000,-336.79,-102.41,-76.094,-40.918,-74.566,-587.69,0.0000,-1054.1,-1530.1,-747.07,-1201.3
1311.000000000,86.215,1868.5,1934.1,1270.8,275.89,2658.4,968.85,1.3463,5442.4,2722.4,3363.4,2052.6,0.0000,-6387.3,-6783.4,-1196.2,-2058.5,-1855.3,-15561.,-105.34,-19201.,-6139.7,-4031.6,-2354.1,61.106,2176.9,1984.9,1300.4,302.75,2762.6,1686.6,0.0000,6478.3,4449.7,4252.8,3658.0,0.0000,-335.22,-101.91,-75.678,-40.737,-73.991,-587.69,0.0000,-1053.9,-1530.0,-747.05,-1201.2
1312.000000000,85.940,1860.5,1925.8,1263.5,274.65,2643.5,968.84,1.3467,5433.7,2722.4,3363.4,2052.8,0.0000,-6381.7,-6780.5,-1194.1,-2057.5,-1851.2,-15559.,-105.30,-19199.,-6139.3,-4031.1,-2353.4,60.836,2167.3,1976.2,1292.7,301.38,2745.4,1686.6,0.0000,6467.9,4449.7,4252.8,3658.0,0.0000,-333.66,-101.41,-75.265,-40.557,-73.417,-587.69,0.0000,-1053.8,-1530.0,-747.04,-1201.1
1313.000000000,85.666,1852.4,1917.4,1256.2,273.36,2628.7,968.84,1.3470,5425.2,2722.4,3363.4,2052.8,0.0000,-6375.9,-6777.6,-1192.0,-2056.5,-1847.0,-15557.,-105.26,-19196.,-6138.9,-4030.6,-2352.7,60.570,2157.8,1967.5,1285.0,300.03,2728.4,1686.6,0.0000,6457.6,4449.7,4252.8,3658.0,0.0000,-332.12,-100.92,-74.855,-40.380,-72.848,-587.69,0.0000,-1053.7,-1529.9,-747.03,-1201.0
1314.000000000,85.396,1844.5,1909.0,1248.9,272.17,2614.1,968.85,1.3474,5417.0,2722.5,3363.4,2052.9,0.0000,-6370.1,-6774.6,-1189.8,-2055.4,-1842.9,-15555.,-105.22,-19194.,-6138.5,-4030.1,-2352.0,60.308,2148.4,1959.0,1277.4,298.69,2711.6,1686.6,0.0000,6447.4,4449.7,4252.8,3658.0,0.0000,-330.60,-100.43,-74.450,-40.205,-72.283,-587.69,0.0000,-1053.6,-1529.8,-747.01,-1200.9
1315.000000000,85.128,1837.0,1900.9,1241.8,271.02,2598.9,968.85,1.3478,5408.2,2722.6,3363.5,2053.0,0.0000,-6364.1,-6771.6,-1187.7,-2054.4,-1838.7,-15553.,-105.18,-19192.,-6138.1,-4029.5,-2351.3,60.050,2139.2,1950.6,1269.8,297.38,2694.9,1686.6,0.0000,6437.4,4449.7,4252.8,3658.0,0.0000,-329.10,-99.947,-74.050,-40.033,-71.723,-587.69,0.0000,-1053.5,-1529.8,-747.00,-1200.8
1316.000000000,84.864,1829.4,1892.8,1234.7,269.88,2583.6,968.85,1.3409,5398.8,2722.6,3363.5,2053.1,0.0000,-6358.1,-6768.6,-1185.5,-2053.3,-1834.4,-15551.,-105.14,-19189.,-6137.7,-4029.0,-2350.6,59.792,2130.1,1942.3,1262.3,296.07,2678.3,1686.6,0.0000,6427.3,4449.7,4252.8,3658.0,0.0000,-327.60,-99.466,-73.651,-39.861,-71.165,-587.69,0.0000,-1053.4,-1529.7,-746.98,-1200.6
1317.000000000,84.601,1821.9,1884.8,1227.6,268.74,2568.2,968.85,1.3372,5389.3,2722.5,3363.5,2053.2,0.0000,-6352.0,-6765.6,-1183.3,-2052.2,-1830.2,-15550.,-105.10,-19187.,-6137.3,-4028.5,-2350.0,59.536,2120.9,1933.9,1254.8,294.76,2661.8,1686.6,0.0000,6417.3,4449.7,4252.8,3658.0,0.0000,-326.11,-98.989,-73.255,-39.691,-70.610,-587.69,0.0000,-1053.3,-1529.6,-746.97,-1200.5
1318.000000000,84.341,1814.3,1876.9,1220.7,267.61,2552.8,968.85,1.3376,5379.8,2722.6,3363.6,2053.3,0.0000,-6345.9,-6762.6,-1181.1,-2051.1,-1825.9,-15548.,-105.06,-19184.,-6136.9,-4028.0,-2349.3,59.284,2112.0,1925.8,1247.4,293.48,2645.4,1686.6,0.0000,6407.4,4449.7,4252.8,3658.0,0.0000,-324.63,-98.517,-72.863,-39.523,-70.060,-587.69,0.0000,-1053.2,-1529.6,-746.96,-1200.4
1319.000000000,84.084,1806.7,1869.2,1213.9,266.49,2537.5,968.85,1.6275,5370.3,2722.6,3363.6,2053.4,0.0000,-6339.8,-6759.6,-1178.9,-2050.1,-1821.6,-15546.,-105.02,-19182.,-6136.5,-4027.5,-2348.6,59.034,2103.1,1917.6,1240.1,292.21,2629.2,1686.6,0.0000,6397.6,4449.7,4252.8,3658.0,0.0000,-323.17,-98.049,-72.474,-39.356,-69.513,-587.69,0.0000,-1053.1,-1529.5,-746.94,-1200.3
1320.000000000,83.829,1800.2,1861.3,1206.8,265.36,2522.3,968.85,2.0010,5361.0,2722.7,3363.6,2053.5,0.0000,-6333.6,-6756.5,-1176.6,-2049.0,-1817.3,-15544.,-104.98,-19179.,-6136.0,-4027.0,-2347.9,58.789,2094.3,1909.7,1232.8,290.96,2613.1,1686.6,0.0000,6387.9,4449.7,4252.8,3658.0,0.0000,-321.74,-97.589,-72.091,-39.192,-68.972,-587.69,0.0000,-1053.0,-1529.4,-746.93,-1200.2
1321.000000000,83.578,1798.3,1858.0,1200.2,264.98,2508.4,968.85,2.0158,5351.8,2722.9,3363.6,2053.6,0.0000,-6327.8,-6753.7,-1174.5,-2047.9,-1813.0,-15542.,-104.95,-19177.,-6135.6,-4026.4,-2347.2,101.78,2137.5,1988.6,1249.0,299.26,2645.7,1686.6,9.8822,6407.4,4451.7,4257.0,3660.7,0.0000,-326.62,-100.10,-73.051,-39.819,-69.659,-587.69,-0.45121,-1053.1,-1529.4,-746.93,-1200.1
1322.000000000,83.855,1810.7,1867.6,1195.7,267.12,2499.3,968.85,2.0162,5343.9,2723.0,3363.6,2053.7,0.0000,-6323.3,-6751.7,-1172.5,-2047.0,-1808.8,-15540.,-104.91,-19174.,-6135.3,-4025.9,-2346.5,250.70,2366.5,2255.8,1282.5,321.66,2700.1,1686.6,603.82,6444.5,4465.2,4271.4,3674.7,0.0000,-334.31,-107.09,-74.450,-40.828,-70.672,-587.69,-27.570,-1053.3,-1529.3,-746.99,-1200.3
1323.000000000,84.605,1833.1,1887.3,1197.3,270.23,2498.8,968.85,2.0165,5337.9,2723.1,3363.6,2053.8,0.0000,-6320.4,-6750.7,-1170.7,-2046.3,-1804.9,-15538.,-104.88,-19172.,-6134.9,-4025.4,-2345.8,72.462,2492.5,2053.5,1359.9,310.69,2836.3,1686.6,58.951,6550.1,4460.0,4253.5,3658.1,0.0000,-338.69,-103.50,-76.284,-41.256,-73.491,-587.69,-2.6916,-1054.2,-1529.2,-746.89,-1199.9
1324.000000000,85.265,1852.9,1906.0,1205.9,273.35,2509.0,968.85,2.0168,5335.9,2723.1,3363.5,2053.9,0.0000,-6318.7,-6750.5,-1169.2,-2045.7,-1801.5,-15536.,-104.84,-19169.,-6134.5,-4024.9,-2345.2,62.283,2218.8,2023.2,1359.2,308.67,2791.5,1686.6,62.475,6543.2,4454.6,4252.9,3658.0,0.0000,-340.59,-103.27,-76.621,-41.524,-73.288,-587.69,-2.8526,-1054.0,-1529.1,-746.87,-1199.8
1325.000000000,86.008,1868.5,1921.2,1218.0,277.03,2522.3,968.86,2.0172,5334.8,2723.2,3363.5,2054.0,0.0000,-6317.7,-6750.6,-1167.8,-2045.2,-1798.5,-15534.,-104.81,-19167.,-6134.1,-4024.3,-2344.5,219.67,2560.2,2385.8,1453.3,363.58,2918.0,1686.6,392.76,6652.6,4506.4,4298.4,3697.3,0.0000,-344.86,-111.67,-77.430,-42.307,-74.377,-587.69,-17.933,-1055.3,-1529.1,-747.09,-1200.4
1326.000000000,86.859,1884.0,1936.3,1228.8,280.06,2534.2,968.81,2.0175,5335.1,2723.3,3363.5,2054.1,0.0000,-6317.5,-6751.1,-1166.6,-2044.7,-1795.9,-15532.,-104.77,-19164.,-6133.7,-4023.8,-2343.8,63.427,2259.5,2060.3,1339.2,316.27,2827.1,1686.6,5.1300,6524.5,4494.6,4273.1,3680.9,0.0000,-346.77,-105.15,-77.841,-42.299,-74.119,-587.69,-0.23423,-1053.4,-1529.0,-746.94,-1200.0
1327.000000000,87.428,1895.8,1948.3,1239.8,281.87,2542.9,968.81,2.4488,5335.0,2723.3,3363.5,2054.2,0.0000,-6317.7,-6751.9,-1165.5,-2044.2,-1793.2,-15530.,-104.73,-19162.,-6133.3,-4023.3,-2343.1,63.432,2259.7,2060.5,1338.0,314.41,2829.0,1686.6,0.0000,6523.9,4459.6,4253.6,3658.4,0.0000,-346.77,-105.15,-77.877,-42.290,-74.137,-587.69,0.0000,-1053.3,-1528.9,-746.83,-1199.5
1328.000000000,87.614,1921.4,1973.0,1254.0,286.19,2567.1,968.81,2.5107,5337.6,2723.4,3363.5,2054.4,0.0000,-6319.1,-6753.4,-1165.2,-2043.9,-1791.0,-15528.,-104.70,-19160.,-6132.9,-4022.8,-2342.5,1187.1,4031.7,3564.9,1735.7,429.65,3563.2,1687.4,2248.1,7037.3,4585.3,4355.1,3753.9,0.0000,-372.83,-141.43,-88.392,-45.718,-90.686,-587.70,-102.65,-1057.0,-1528.9,-747.33,-1201.1
1329.000000000,90.135,1981.9,2026.3,1293.9,295.87,2643.4,968.81,2.5110,5360.3,2723.4,3363.7,2054.5,0.0000,-6324.0,-6757.0,-1166.1,-2044.0,-1790.2,-15526.,-104.67,-19158.,-6132.5,-4022.2,-2341.8,69.174,2606.0,2256.9,1983.1,451.28,3662.1,1686.6,270.44,7249.4,4772.0,4530.0,3956.9,0.0000,-378.44,-114.97,-89.641,-46.772,-91.596,-587.69,-12.348,-1059.9,-1528.8,-748.19,-1204.6
1330.000000000,91.543,2029.8,2075.5,1357.3,304.37,2737.0,968.81,2.5114,5391.1,2723.5,3364.4,2054.9,0.0000,-6331.0,-6761.9,-1166.8,-2044.2,-1791.2,-15524.,-104.63,-19156.,-6132.1,-4021.7,-2341.1,69.752,2811.2,2368.8,1913.0,432.18,3744.0,1694.3,457.24,7205.6,4743.9,4530.7,3938.0,0.0000,-381.95,-117.98,-90.561,-47.021,-92.865,-587.80,-20.877,-1059.0,-1528.7,-748.18,-1204.1
1331.000000000,92.590,2057.4,2104.5,1401.6,310.50,2816.2,968.78,33.072,5430.5,2724.2,3366.4,2055.9,0.0000,-6338.3,-6766.8,-1168.2,-2044.5,-1793.3,-15522.,-104.60,-19154.,-6131.7,-4021.2,-2340.4,252.49,2672.2,2419.9,1908.1,475.23,3780.2,1702.3,623.37,7212.6,4718.5,4511.5,3918.2,0.0000,-384.29,-119.59,-91.513,-47.577,-94.136,-587.92,-28.462,-1058.7,-1528.7,-748.07,-1203.7
1332.000000000,93.926,2075.0,2126.0,1451.5,313.99,2882.0,968.78,42.058,5463.7,2731.7,3369.2,2058.8,0.0000,-6345.6,-6771.5,-1169.6,-2044.6,-1794.8,-15520.,-104.57,-19153.,-6131.4,-4020.7,-2339.8,70.371,2506.9,2285.9,1694.2,377.78,3597.0,1686.6,0.0000,7005.7,4498.2,4296.8,3702.2,0.0000,-384.98,-116.95,-92.021,-47.078,-94.005,-587.69,0.0000,-1055.6,-1528.6,-746.98,-1199.7
1333.000000000,94.380,2087.3,2138.1,1481.8,315.35,2939.5,968.78,32.478,5493.4,2737.8,3375.7,2061.1,0.0000,-6352.4,-6775.7,-1171.4,-2044.7,-1795.8,-15518.,-104.53,-19151.,-6131.1,-4020.2,-2339.1,70.269,2503.3,2282.6,1676.9,359.94,3600.4,1686.6,0.0000,6995.4,4469.6,4271.0,3676.3,0.0000,-384.51,-116.85,-92.308,-46.902,-94.630,-587.69,0.0000,-1055.2,-1528.6,-746.84,-1199.2
1334.000000000,94.510,2092.2,2143.5,1510.6,315.70,2978.5,968.78,50.308,5528.4,2746.0,3371.5,2062.6,0.0000,-6358.5,-6779.4,-1173.6,-2044.7,-1796.7,-15516.,-104.50,-19149.,-6131.0,-4019.7,-2338.4,70.061,2495.9,2275.8,1669.1,353.64,3610.5,1686.6,0.0000,6994.5,4459.6,4264.4,3672.3,0.0000,-383.45,-116.57,-92.452,-46.729,-95.160,-587.69,0.0000,-1055.0,-1528.5,-746.79,-1199.0
1335.000000000,94.468,2091.6,2146.0,1528.3,315.39,3019.6,968.75,65.058,5577.8,2738.2,3371.0,2061.7,0.0000,-6363.8,-6782.5,-1175.4,-2044.6,-1797.3,-15514.,-104.46,-19148.,-6131.0,-4019.2,-2337.8,69.806,2486.8,2267.5,1670.0,349.34,3623.6,1686.6,0.0000,7000.4,4451.5,4255.1,3661.2,0.0000,-382.13,-116.20,-92.528,-46.539,-95.640,-587.69,0.0000,-1055.0,-1528.4,-746.74,-1198.7
1336.000000000,94.296,2092.0,2147.4,1539.2,314.71,3085.2,968.75,71.639,5642.5,2733.6,3369.1,2060.6,0.0000,-6368.5,-6785.2,-1176.9,-2044.4,-1797.8,-15512.,-104.43,-19147.,-6130.9,-4018.7,-2337.1,69.587,2479.0,2260.4,1674.5,348.08,3638.7,1686.6,0.0000,7009.3,4449.7,4252.9,3658.2,0.0000,-381.00,-115.89,-92.599,-46.391,-96.078,-587.69,0.0000,-1055.0,-1528.4,-746.72,-1198.6
1337.000000000,94.147,2090.5,2146.2,1548.0,313.98,3151.5,968.75,66.189,5688.6,2731.7,3367.3,2061.1,0.0000,-6372.6,-6787.5,-1178.2,-2044.1,-1798.3,-15510.,-104.39,-19146.,-6130.8,-4018.3,-2336.5,69.410,2472.7,2254.7,1680.3,347.37,3655.8,1686.6,125.40,7019.8,4557.9,4252.8,3670.6,0.0000,-380.10,-115.63,-92.715,-46.273,-96.557,-587.69,-5.7255,-1055.0,-1528.3,-746.71,-1198.7
1338.000000000,94.068,2087.3,2143.2,1558.1,313.26,3197.3,968.75,47.561,5721.0,2729.7,3367.1,2061.0,0.0000,-6376.2,-6789.4,-1179.4,-2043.8,-1798.7,-15508.,-104.36,-19145.,-6130.5,-4017.8,-2335.9,69.227,2466.2,2248.7,1684.8,346.61,3669.5,1686.6,0.0000,7028.1,4449.7,4252.8,3658.0,0.0000,-379.15,-115.36,-92.781,-46.151,-96.942,-587.69,0.0000,-1055.0,-1528.2,-746.71,-1198.4
1339.000000000,93.866,2086.4,2139.7,1570.7,312.55,3226.1,968.75,54.001,5743.8,2732.0,3366.3,2060.4,0.0000,-6379.0,-6791.1,-1180.6,-2043.5,-1799.1,-15507.,-104.32,-19144.,-6130.3,-4017.3,-2335.2,68.987,2457.6,2240.9,1688.8,345.57,3682.6,1686.6,123.45,7036.1,4474.5,4252.8,3658.0,0.0000,-377.89,-115.00,-92.802,-45.991,-97.313,-587.69,-5.6365,-1055.0,-1528.2,-746.70,-1198.3
1340.000000000,93.646,2082.8,2136.9,1579.3,311.92,3245.9,968.71,51.668,5760.6,2733.1,3365.9,2060.1,0.0000,-6381.3,-6792.5,-1181.6,-2043.2,-1799.6,-15505.,-104.29,-19143.,-6130.1,-4016.8,-2334.6,68.694,2447.2,2231.4,1691.3,344.27,3692.5,1686.6,0.0000,7042.2,4449.7,4252.8,3658.0,0.0000,-376.33,-114.54,-92.746,-45.796,-97.598,-587.69,0.0000,-1055.0,-1528.1,-746.69,-1198.2
1341.000000000,93.607,2076.7,2131.5,1584.7,311.09,3262.6,968.71,43.217,5770.2,2735.0,3365.9,2059.6,0.0000,-6383.0,-6793.7,-1182.6,-2042.8,-1800.1,-15503.,-104.25,-19142.,-6129.8,-4016.4,-2333.9,68.464,2439.0,2223.9,1693.0,343.24,3699.5,1686.6,0.0000,7046.5,4449.7,4252.8,3658.0,0.0000,-375.10,-114.18,-92.692,-45.642,-97.801,-587.69,0.0000,-1055.0,-1528.1,-746.68,-1198.1
1342.000000000,93.405,2072.3,2126.2,1589.0,310.14,3280.4,968.71,38.238,5779.3,2734.1,3366.5,2059.7,0.0000,-6384.3,-6794.6,-1183.5,-2042.4,-1800.6,-15501.,-104.21,-19141.,-6129.6,-4015.9,-2333.3,68.228,2430.6,2216.3,1764.6,342.21,3709.5,1686.6,413.28,7253.7,4654.8,4394.9,3859.0,0.0000,-373.84,-113.80,-92.675,-45.485,-98.089,-587.69,-18.870,-1057.8,-1528.0,-747.38,-1201.5
1343.000000000,93.154,2065.9,2121.7,1592.3,309.13,3298.4,968.72,31.089,5793.9,2732.8,3366.4,2059.5,0.0000,-6385.3,-6795.3,-1184.4,-2042.0,-1801.3,-15500.,-104.18,-19140.,-6129.3,-4015.4,-2332.6,67.910,2419.3,2206.0,1695.0,340.74,3710.8,1686.6,0.0000,7053.5,4449.7,4252.8,3658.0,0.0000,-372.12,-113.28,-92.488,-45.273,-98.139,-587.69,0.0000,-1054.9,-1527.9,-746.66,-1197.9
1344.000000000,92.866,2059.1,2114.0,1595.3,308.01,3319.0,968.72,26.989,5805.3,2732.2,3365.9,2060.3,0.0000,-6385.9,-6795.6,-1185.1,-2041.5,-1802.0,-15498.,-104.14,-19139.,-6129.0,-4014.9,-2332.0,67.578,2407.4,2195.2,1693.3,339.18,3710.4,1686.6,0.0000,7053.3,4449.7,4252.8,3658.0,0.0000,-370.32,-112.74,-92.269,-45.052,-98.142,-587.69,0.0000,-1054.9,-1527.9,-746.64,-1197.8
1345.000000000,92.638,2050.8,2105.4,1600.1,306.78,3330.1,968.72,26.311,5811.6,2731.8,3365.7,2061.1,0.0000,-6385.9,-6795.6,-1185.8,-2040.9,-1802.7,-15496.,-104.11,-19138.,-6128.8,-4014.4,-2331.3,67.249,2395.7,2184.5,1691.2,337.64,3708.5,1686.6,0.0000,7052.2,4449.7,4252.8,3658.0,0.0000,-368.53,-112.19,-92.033,-44.833,-98.105,-587.69,0.0000,-1054.9,-1527.8,-746.63,-1197.7
1346.000000000,92.361,2041.8,2096.7,1600.6,305.49,3338.4,968.72,26.319,5818.1,2733.9,3365.7,2061.1,0.0000,-6385.5,-6795.4,-1186.4,-2040.4,-1803.4,-15494.,-104.07,-19138.,-6128.5,-4013.9,-2330.7,66.920,2384.0,2173.8,1688.5,336.08,3705.2,1686.6,0.0000,7050.3,4449.7,4252.8,3658.0,0.0000,-366.73,-111.64,-91.777,-44.613,-98.026,-587.69,0.0000,-1054.8,-1527.7,-746.62,-1197.6
1347.000000000,92.031,2032.8,2088.6,1600.8,304.14,3342.0,968.72,22.916,5827.2,2733.2,3365.7,2061.3,0.0000,-6384.6,-6794.9,-1186.9,-2039.8,-1804.0,-15493.,-104.03,-19137.,-6128.2,-4013.4,-2330.0,66.593,2372.4,2163.2,1685.3,334.53,3700.6,1686.6,0.0000,7047.5,4449.7,4252.8,3658.0,0.0000,-364.94,-111.09,-91.505,-44.396,-97.911,-587.69,0.0000,-1054.8,-1527.7,-746.61,-1197.5
1348.000000000,91.701,2024.4,2079.9,1600.0,302.82,3346.7,968.72,20.760,5832.3,2734.7,3365.6,2061.4,0.0000,-6383.4,-6794.1,-1187.3,-2039.1,-1804.6,-15491.,-104.00,-19136.,-6128.0,-4012.9,-2329.4,66.270,2360.8,2152.7,1681.7,332.98,3694.8,1686.6,0.0000,7044.1,4449.7,4252.8,3658.0,0.0000,-363.16,-110.54,-91.220,-44.180,-97.763,-587.69,0.0000,-1054.7,-1527.6,-746.59,-1197.4
1349.000000000,91.525,2016.2,2071.0,1598.2,301.49,3352.0,968.72,16.771,5839.3,2734.7,3365.6,2061.6,0.0000,-6381.8,-6793.1,-1187.6,-2038.5,-1805.2,-15489.,-103.96,-19135.,-6127.7,-4012.4,-2328.7,65.956,2349.6,2142.5,1677.8,331.47,3688.3,1686.6,0.0000,7040.2,4449.7,4252.8,3658.0,0.0000,-361.42,-110.00,-90.931,-43.971,-97.594,-587.69,0.0000,-1054.7,-1527.5,-746.58,-1197.3
1350.000000000,90.980,2008.2,2063.5,1596.8,300.33,3351.9,968.70,16.770,5842.5,2733.7,3366.0,2061.9,0.0000,-6380.0,-6791.9,-1187.9,-2037.8,-1805.8,-15488.,-103.92,-19134.,-6127.5,-4011.9,-2328.1,65.829,2356.8,2138.4,1676.6,330.87,3686.5,1686.6,0.0000,7039.1,4449.7,4252.8,3658.0,0.0000,-360.72,-109.77,-90.826,-43.886,-97.550,-587.69,0.0000,-1054.6,-1527.5,-746.56,-1197.2
1351.000000000,90.341,2001.6,2058.2,1594.8,299.37,3354.6,968.70,16.769,5845.6,2733.6,3366.4,2061.8,0.0000,-6378.0,-6790.7,-1188.1,-2037.1,-1806.3,-15486.,-103.89,-19134.,-6127.2,-4011.4,-2327.4,65.534,2334.6,2128.8,1672.2,329.44,3678.5,1686.6,0.0000,7034.3,4449.7,4252.8,3658.0,0.0000,-359.07,-109.26,-90.529,-43.690,-97.335,-587.69,0.0000,-1054.6,-1527.4,-746.55,-1197.1
1352.000000000,89.867,1995.0,2055.8,1592.8,298.38,3358.2,968.68,14.178,5850.5,2734.9,3366.1,2061.7,0.0000,-6376.1,-6789.4,-1188.2,-2036.4,-1806.7,-15485.,-103.85,-19133.,-6127.0,-4010.9,-2326.8,65.470,2352.6,2127.6,1684.5,329.15,3679.1,1686.6,60.078,7049.8,4535.7,4318.8,3778.0,0.0000,-358.72,-109.15,-90.497,-43.647,-97.353,-587.69,-2.7431,-1054.8,-1527.4,-746.87,-1199.1
1353.000000000,89.681,1990.0,2051.1,1590.6,297.80,3357.0,968.66,14.393,5858.5,2733.1,3365.8,2061.4,0.0000,-6374.1,-6788.1,-1188.3,-2035.7,-1807.0,-15483.,-103.81,-19132.,-6126.7,-4010.4,-2326.1,65.218,2323.4,2118.5,1668.1,327.92,3671.4,1686.6,0.0000,7030.1,4449.7,4252.8,3658.0,0.0000,-357.28,-108.69,-90.231,-43.479,-97.146,-587.69,0.0000,-1054.5,-1527.3,-746.52,-1196.9
1354.000000000,89.468,1983.6,2045.7,1588.4,296.84,3356.7,968.66,14.533,5860.4,2733.0,3365.6,2061.2,0.0000,-6372.0,-6786.7,-1188.3,-2035.0,-1807.3,-15482.,-103.78,-19131.,-6126.4,-4009.9,-2325.5,65.006,2315.8,2111.6,1664.8,326.89,3665.2,1686.6,0.0000,7026.4,4449.7,4252.8,3658.0,0.0000,-356.08,-108.31,-90.012,-43.337,-96.978,-587.69,0.0000,-1054.4,-1527.2,-746.51,-1196.8
1355.000000000,89.258,1976.6,2040.3,1586.5,295.99,3357.9,968.66,16.793,5861.4,2733.6,3366.0,2061.3,0.0000,-6369.8,-6785.1,-1188.3,-2034.2,-1807.6,-15480.,-103.74,-19130.,-6126.1,-4009.4,-2324.8,64.721,2305.7,2102.4,1659.1,325.49,3653.8,1686.6,0.0000,7019.5,4449.7,4252.8,3658.0,0.0000,-354.49,-107.81,-89.674,-43.147,-96.666,-587.69,0.0000,-1054.4,-1527.2,-746.50,-1196.7
1356.000000000,88.970,1968.9,2034.5,1583.4,294.88,3356.9,968.66,15.747,5861.8,2733.8,3366.1,2061.6,0.0000,-6367.4,-6783.4,-1188.2,-2033.5,-1808.1,-15479.,-103.70,-19129.,-6125.8,-4008.9,-2324.2,64.438,2295.6,2093.2,1653.2,324.09,3641.6,1686.6,0.0000,7012.1,4449.7,4252.8,3658.0,0.0000,-352.90,-107.31,-89.329,-42.959,-96.332,-587.69,0.0000,-1054.3,-1527.1,-746.48,-1196.6
1357.000000000,88.792,1960.6,2027.0,1579.3,293.75,3352.8,968.66,13.642,5859.7,2733.9,3366.0,2061.5,0.0000,-6364.8,-6781.6,-1188.1,-2032.7,-1808.5,-15477.,-103.67,-19128.,-6125.5,-4008.4,-2323.5,64.156,2285.5,2084.0,1647.1,322.68,3628.7,1686.6,0.0000,7004.4,4449.7,4252.8,3658.0,0.0000,-351.31,-106.81,-88.973,-42.770,-95.977,-587.69,0.0000,-1054.3,-1527.0,-746.47,-1196.5
1358.000000000,88.575,1952.8,2019.3,1574.7,292.57,3347.5,968.66,14.392,5856.9,2734.7,3365.6,2061.2,0.0000,-6361.9,-6779.6,-1187.9,-2031.9,-1808.7,-15476.,-103.63,-19127.,-6125.2,-4007.9,-2322.8,63.873,2275.4,2074.8,1640.6,321.28,3615.1,1686.6,0.0000,6996.1,4449.7,4252.8,3658.0,0.0000,-349.71,-106.31,-88.608,-42.582,-95.601,-587.69,0.0000,-1054.2,-1527.0,-746.45,-1196.4
1359.000000000,88.126,1944.6,2011.2,1569.6,291.36,3344.1,968.66,13.744,5854.3,2734.6,3365.6,2061.2,0.0000,-6358.8,-6777.5,-1187.5,-2031.1,-1808.6,-15474.,-103.59,-19126.,-6124.9,-4007.4,-2322.2,63.593,2265.5,2065.7,1634.0,319.88,3601.1,1686.6,0.0000,6987.6,4449.7,4252.8,3658.0,0.0000,-348.13,-105.81,-88.237,-42.395,-95.210,-587.69,0.0000,-1054.1,-1526.9,-746.44,-1196.3
1360.000000000,87.852,1936.8,2003.1,1564.1,290.15,3338.0,968.67,14.011,5850.6,2735.1,3365.5,2061.4,0.0000,-6355.4,-6775.4,-1187.2,-2030.2,-1808.4,-15473.,-103.56,-19125.,-6124.6,-4006.9,-2321.5,63.326,2255.9,2057.0,1627.4,318.54,3586.9,1686.6,0.0000,6979.1,4449.7,4252.8,3658.0,0.0000,-346.61,-105.33,-87.874,-42.217,-94.815,-587.69,0.0000,-1054.1,-1526.8,-746.43,-1196.2
1361.000000000,87.514,1929.0,1994.9,1558.4,288.97,3333.0,968.67,15.293,5846.2,2734.0,3365.4,2061.5,0.0000,-6351.9,-6773.2,-1186.7,-2029.4,-1808.1,-15471.,-103.52,-19124.,-6124.2,-4006.4,-2320.9,63.066,2246.7,2048.6,1620.7,317.23,3572.5,1686.6,0.0000,6970.4,4449.7,4252.8,3658.0,0.0000,-345.13,-104.86,-87.511,-42.044,-94.410,-587.69,0.0000,-1054.0,-1526.8,-746.41,-1196.1
1362.000000000,87.036,1921.0,1987.0,1552.6,287.82,3324.4,968.67,15.297,5841.4,2733.5,3365.3,2062.0,0.0000,-6348.2,-6770.9,-1186.2,-2028.5,-1807.6,-15470.,-103.48,-19123.,-6123.9,-4005.9,-2320.2,62.809,2237.5,2040.3,1613.8,315.93,3557.6,1686.6,0.0000,6961.4,4449.7,4252.8,3658.0,0.0000,-343.67,-104.40,-87.144,-41.873,-93.991,-587.69,0.0000,-1053.9,-1526.7,-746.40,-1196.0
1363.000000000,86.704,1913.3,1979.0,1546.5,286.68,3318.0,968.64,13.661,5836.5,2733.5,3365.2,2062.3,0.0000,-6344.3,-6768.6,-1185.6,-2027.6,-1807.0,-15468.,-103.44,-19123.,-6123.6,-4005.5,-2319.6,62.553,2228.4,2031.9,1606.8,314.64,3542.3,1686.6,0.0000,6952.1,4449.7,4252.8,3658.0,0.0000,-342.20,-103.93,-86.772,-41.702,-93.559,-587.69,0.0000,-1053.8,-1526.6,-746.38,-1195.9
1364.000000000,86.587,1917.8,1982.3,1541.1,287.60,3309.6,968.63,13.035,5834.9,2733.5,3365.2,2062.5,0.0000,-6341.1,-6766.8,-1185.2,-2026.8,-1806.3,-15467.,-103.41,-19122.,-6123.3,-4005.0,-2318.9,120.28,2410.9,2170.2,1663.1,335.46,3611.9,1686.6,134.94,7012.4,4488.1,4281.0,3694.8,0.0000,-355.89,-109.26,-89.116,-43.412,-95.047,-587.69,-6.1612,-1054.3,-1526.6,-746.51,-1196.4
1365.000000000,87.822,1990.1,2045.9,1551.0,299.98,3345.3,968.60,13.145,5837.3,2733.3,3365.5,2061.9,0.0000,-6343.0,-6768.4,-1186.3,-2026.7,-1806.8,-15465.,-103.38,-19122.,-6122.9,-4004.5,-2318.3,2696.9,5275.8,4701.9,2065.6,408.28,4482.5,1691.7,2167.5,7560.5,4531.3,4318.7,3737.1,0.0000,-412.46,-172.64,-106.48,-49.953,-117.94,-587.76,-98.965,-1056.9,-1526.5,-746.68,-1197.0
1366.000000000,93.547,2162.8,2197.5,1623.3,327.32,3481.0,968.60,11.387,5869.4,2733.9,3366.1,2061.5,0.0000,-6355.8,-6777.0,-1188.7,-2027.9,-1810.1,-15464.,-103.35,-19121.,-6122.6,-4004.0,-2317.6,191.26,3046.9,2817.6,2655.8,718.09,4862.7,1706.3,175.84,8149.6,5099.4,4780.9,4240.0,0.0000,-451.20,-140.16,-111.84,-56.819,-119.97,-587.97,-8.0285,-1065.2,-1526.4,-748.98,-1205.6
1367.000000000,99.444,2319.7,2351.1,1720.6,350.82,3619.3,968.59,11.387,5912.9,2734.5,3368.1,2063.1,0.0000,-6376.5,-6790.7,-1191.8,-2029.9,-1816.6,-15462.,-103.32,-19121.,-6122.3,-4003.5,-2317.0,83.083,2959.8,2698.8,2091.5,469.64,4511.4,1689.9,0.0000,7548.9,4518.3,4322.1,3736.2,0.0000,-454.97,-138.51,-112.32,-55.717,-118.51,-587.74,0.0000,-1056.7,-1526.4,-746.67,-1196.8
1368.000000000,103.14,2387.5,2427.7,1798.8,366.15,3699.2,968.55,19.209,5943.3,2741.5,3368.5,2065.6,0.0000,-6398.3,-6804.0,-1195.3,-2031.7,-1822.4,-15461.,-103.29,-19121.,-6121.9,-4003.0,-2316.3,83.040,2958.3,2697.5,2075.6,446.86,4486.1,1689.5,0.0000,7531.9,4492.8,4294.2,3704.6,0.0000,-455.01,-138.66,-112.29,-55.549,-118.46,-587.73,0.0000,-1056.4,-1526.3,-746.52,-1196.2
1369.000000000,107.05,2412.4,2461.0,1845.8,372.97,3750.9,968.56,31.453,5969.1,2744.3,3371.6,2066.3,0.0000,-6419.3,-6815.1,-1199.3,-2033.2,-1826.9,-15459.,-103.26,-19121.,-6121.7,-4002.6,-2315.7,82.812,2950.1,2690.0,2054.6,426.55,4461.9,1689.5,0.0000,7510.6,4466.5,4268.9,3676.6,0.0000,-454.06,-138.49,-112.12,-55.279,-118.38,-587.73,0.0000,-1056.2,-1526.3,-746.38,-1195.6
1370.000000000,108.14,2422.8,2475.4,1872.4,372.72,3775.7,968.56,39.505,6013.0,2745.1,3369.5,2067.5,0.0000,-6438.0,-6824.8,-1203.6,-2034.2,-1830.6,-15458.,-103.22,-19121.,-6121.5,-4002.1,-2315.0,82.494,2938.8,2679.7,2043.5,416.92,4447.9,1689.2,0.0000,7499.5,4455.1,4258.0,3664.3,0.0000,-452.61,-138.17,-111.87,-55.017,-118.31,-587.73,0.0000,-1056.0,-1526.2,-746.32,-1195.3
1371.000000000,107.90,2427.6,2482.1,1882.4,371.54,3823.9,968.56,27.170,6098.8,2740.5,3369.9,2066.9,0.0000,-6455.0,-6833.3,-1206.9,-2035.0,-1833.8,-15456.,-103.19,-19121.,-6121.4,-4001.6,-2314.4,82.129,2925.8,2667.9,2036.8,412.27,4438.1,1689.0,0.0000,7492.9,4450.6,4253.7,3659.2,0.0000,-450.90,-137.75,-111.57,-54.756,-118.21,-587.72,0.0000,-1056.0,-1526.2,-746.28,-1195.1
1372.000000000,107.54,2425.9,2493.6,1881.5,370.10,3914.5,968.56,38.045,6177.1,2738.3,3369.1,2067.6,0.0000,-6470.9,-6840.5,-1209.6,-2035.7,-1836.6,-15455.,-103.15,-19120.,-6121.1,-4001.2,-2313.8,81.735,2911.8,2655.1,2031.6,409.96,4429.5,1689.0,0.0000,7487.7,4449.7,4252.8,3658.0,0.0000,-449.00,-137.26,-111.22,-54.490,-118.08,-587.72,0.0000,-1056.0,-1526.1,-746.27,-1195.0
1373.000000000,106.49,2432.9,2500.9,1880.8,368.49,3981.0,968.56,41.125,6223.2,2738.6,3368.4,2067.7,0.0000,-6485.9,-6847.0,-1211.8,-2036.1,-1839.0,-15454.,-103.12,-19121.,-6120.9,-4000.8,-2313.2,81.323,2897.1,2641.7,2026.2,407.98,4420.1,1688.8,0.0000,7482.1,4449.7,4252.8,3658.0,0.0000,-446.99,-136.72,-110.84,-54.216,-117.91,-587.72,0.0000,-1055.9,-1526.0,-746.26,-1194.9
1374.000000000,105.96,2426.1,2490.6,1896.3,366.76,3992.4,968.56,33.058,6240.1,2740.9,3367.9,2066.9,0.0000,-6499.1,-6852.4,-1213.9,-2036.5,-1841.3,-15452.,-103.08,-19121.,-6120.6,-4000.3,-2312.5,80.888,2881.6,2627.5,2020.0,405.87,4408.9,1688.6,0.0000,7475.3,4449.7,4252.8,3658.0,0.0000,-444.83,-136.12,-110.43,-53.925,-117.69,-587.72,0.0000,-1055.9,-1526.0,-746.25,-1194.8
1375.000000000,105.39,2422.4,2478.3,1903.0,364.97,3987.6,968.57,34.148,6244.4,2740.7,3367.8,2066.7,0.0000,-6510.3,-6857.2,-1215.8,-2036.8,-1843.4,-15451.,-103.05,-19121.,-6120.4,-3999.9,-2311.9,80.448,2865.9,2613.2,2013.3,403.74,4396.6,1688.6,0.0000,7467.9,4449.7,4252.8,3658.0,0.0000,-442.62,-135.50,-109.99,-53.632,-117.43,-587.72,0.0000,-1055.9,-1525.9,-746.24,-1194.7
1376.000000000,104.96,2420.5,2474.1,1899.2,363.17,3983.0,968.57,35.550,6240.5,2739.9,3367.3,2066.5,0.0000,-6519.9,-6861.5,-1217.5,-2037.0,-1845.4,-15450.,-103.01,-19121.,-6120.1,-3999.4,-2311.3,80.011,2850.3,2599.0,2006.4,401.61,4383.5,1688.5,0.0000,7460.1,4449.7,4252.8,3658.0,0.0000,-440.41,-134.88,-109.54,-53.340,-117.15,-587.71,0.0000,-1055.8,-1525.9,-746.23,-1194.6
1377.000000000,104.52,2409.9,2467.3,1893.8,361.55,3988.0,968.57,33.792,6241.7,2739.5,3367.1,2066.6,0.0000,-6528.1,-6865.2,-1219.0,-2037.2,-1847.4,-15448.,-102.98,-19121.,-6119.8,-3999.0,-2310.7,79.616,2836.3,2586.2,2000.2,399.70,4371.8,1688.3,0.0000,7453.1,4449.7,4252.8,3658.0,0.0000,-438.41,-134.31,-109.14,-53.077,-116.90,-587.71,0.0000,-1055.8,-1525.8,-746.22,-1194.6
1378.000000000,104.09,2403.8,2457.7,1888.1,359.78,3995.2,968.57,30.454,6247.8,2738.6,3367.8,2067.8,0.0000,-6535.4,-6868.7,-1220.4,-2037.3,-1849.4,-15447.,-102.94,-19121.,-6119.5,-3998.5,-2310.1,79.218,2822.1,2573.3,1993.4,397.75,4358.7,1688.2,0.0000,7445.2,4449.7,4252.8,3658.0,0.0000,-436.38,-133.73,-108.72,-52.812,-116.60,-587.71,0.0000,-1055.8,-1525.8,-746.21,-1194.5
1379.000000000,103.46,2392.8,2458.9,1888.0,358.08,3994.3,968.57,29.399,6242.9,2738.0,3367.4,2067.8,0.0000,-6542.8,-6871.7,-1221.6,-2037.3,-1851.4,-15446.,-102.91,-19121.,-6119.3,-3998.1,-2309.5,78.830,2808.3,2560.7,1986.5,395.85,4345.1,1687.1,0.0000,7437.0,4449.7,4252.8,3658.0,0.0000,-434.39,-133.15,-108.29,-52.554,-116.31,-587.70,0.0000,-1055.7,-1525.7,-746.20,-1194.4
1380.000000000,102.94,2384.6,2447.1,1884.8,356.39,3987.7,968.57,26.677,6239.2,2737.9,3366.9,2067.2,0.0000,-6549.2,-6874.2,-1222.7,-2037.3,-1853.3,-15444.,-102.87,-19121.,-6119.0,-3997.6,-2308.8,78.445,2794.6,2548.2,1979.3,393.96,4330.8,1686.8,0.0000,7428.4,4449.7,4252.8,3658.0,0.0000,-432.40,-132.56,-107.86,-52.297,-115.99,-587.69,0.0000,-1055.7,-1525.6,-746.19,-1194.3
1381.000000000,102.46,2376.6,2435.7,1879.3,354.68,3976.2,968.58,22.786,6241.1,2738.7,3366.8,2067.2,0.0000,-6554.7,-6876.4,-1223.6,-2037.2,-1855.1,-15443.,-102.84,-19121.,-6118.7,-3997.2,-2308.2,78.057,2780.7,2535.6,1971.8,392.05,4315.6,1686.7,0.0000,7419.2,4449.7,4252.8,3658.0,0.0000,-430.38,-131.97,-107.41,-52.038,-115.65,-587.69,0.0000,-1055.6,-1525.6,-746.18,-1194.2
1382.000000000,102.16,2365.0,2424.0,1873.0,353.01,3970.9,968.58,20.722,6237.9,2738.7,3366.6,2066.9,0.0000,-6559.3,-6878.2,-1224.5,-2037.1,-1856.9,-15442.,-102.80,-19121.,-6118.4,-3996.7,-2307.6,77.662,2766.7,2522.7,1963.8,390.10,4299.3,1686.6,0.0000,7409.4,4449.7,4252.8,3658.0,0.0000,-428.32,-131.35,-106.94,-51.775,-115.28,-587.69,0.0000,-1055.6,-1525.5,-746.17,-1194.1
1383.000000000,101.75,2353.0,2412.7,1868.6,351.30,3961.7,968.58,18.888,6234.1,2737.7,3366.5,2066.5,0.0000,-6563.2,-6879.6,-1225.2,-2036.9,-1858.6,-15441.,-102.76,-19120.,-6118.1,-3996.3,-2306.9,77.277,2752.9,2510.2,1955.7,388.20,4282.7,1686.6,0.0000,7399.3,4449.7,4252.8,3658.0,0.0000,-426.29,-130.74,-106.48,-51.518,-114.89,-587.69,0.0000,-1055.6,-1525.5,-746.16,-1194.0
1384.000000000,101.36,2341.8,2400.8,1862.7,349.63,3954.3,968.58,18.574,6229.7,2737.5,3366.7,2066.3,0.0000,-6566.2,-6880.5,-1225.8,-2036.6,-1860.2,-15439.,-102.73,-19120.,-6117.8,-3995.8,-2306.3,76.887,2739.0,2497.6,1947.3,386.26,4265.2,1686.6,0.0000,7388.8,4449.7,4252.8,3658.0,0.0000,-424.22,-130.11,-105.99,-51.258,-114.47,-587.69,0.0000,-1055.5,-1525.4,-746.14,-1193.9
1385.000000000,100.97,2332.6,2389.3,1856.9,347.93,3948.1,968.58,16.628,6229.9,2738.0,3366.5,2066.6,0.0000,-6568.6,-6881.0,-1226.3,-2036.3,-1861.6,-15438.,-102.69,-19120.,-6117.5,-3995.4,-2305.7,76.496,2725.1,2484.9,1938.6,384.32,4247.0,1686.6,0.0000,7377.8,4449.7,4252.8,3658.0,0.0000,-422.13,-129.47,-105.50,-50.997,-114.02,-587.69,0.0000,-1055.4,-1525.3,-746.13,-1193.8
1386.000000000,100.57,2320.9,2380.1,1851.4,346.25,3933.7,968.58,16.628,6233.8,2737.9,3366.7,2066.3,0.0000,-6570.3,-6881.1,-1226.7,-2036.0,-1862.7,-15437.,-102.66,-19119.,-6117.1,-3994.9,-2305.0,76.109,2711.3,2472.3,1929.7,382.39,4228.3,1686.6,0.0000,7366.5,4449.7,4252.8,3658.0,0.0000,-420.05,-128.83,-105.00,-50.739,-113.56,-587.69,0.0000,-1055.4,-1525.3,-746.12,-1193.7
1387.000000000,100.18,2309.2,2374.7,1843.8,344.57,3924.9,968.57,14.706,6227.2,2737.2,3367.0,2066.0,0.0000,-6571.7,-6881.0,-1227.0,-2035.6,-1863.7,-15436.,-102.62,-19119.,-6116.8,-3994.5,-2304.4,75.728,2697.8,2459.9,1920.8,380.49,4209.4,1686.6,0.0000,7355.1,4449.7,4252.8,3658.0,0.0000,-418.00,-128.19,-104.50,-50.486,-113.09,-587.69,0.0000,-1055.3,-1525.2,-746.10,-1193.6
1388.000000000,99.798,2300.5,2372.2,1835.9,342.89,3915.0,968.54,14.620,6223.9,2736.5,3366.9,2066.0,0.0000,-6573.0,-6880.6,-1227.2,-2035.2,-1864.9,-15435.,-102.58,-19119.,-6116.4,-3994.0,-2303.7,75.353,2684.4,2447.7,1911.7,378.61,4190.1,1686.6,0.0000,7343.4,4449.7,4252.8,3658.0,0.0000,-415.97,-127.56,-104.01,-50.235,-112.60,-587.69,0.0000,-1055.3,-1525.2,-746.09,-1193.5
1389.000000000,99.387,2289.7,2360.5,1827.8,341.26,3902.2,968.54,12.787,6215.3,2736.0,3367.2,2065.7,0.0000,-6573.9,-6879.9,-1227.3,-2034.8,-1866.1,-15434.,-102.55,-19118.,-6116.1,-3993.6,-2303.1,74.995,2671.7,2436.1,1902.9,376.82,4171.0,1686.6,0.0000,7331.9,4449.7,4252.8,3658.0,0.0000,-414.02,-126.95,-103.52,-49.997,-112.12,-587.69,0.0000,-1055.2,-1525.1,-746.08,-1193.4
1390.000000000,98.953,2279.0,2349.8,1821.4,339.67,3888.2,968.54,12.623,6208.7,2735.6,3367.2,2065.6,0.0000,-6574.3,-6878.9,-1227.3,-2034.3,-1867.1,-15432.,-102.51,-19118.,-6115.7,-3993.1,-2302.4,74.680,2660.4,2425.9,1894.8,375.23,4153.7,1686.6,0.0000,7321.4,4449.7,4252.8,3658.0,0.0000,-412.30,-126.41,-103.08,-49.787,-111.67,-587.69,0.0000,-1055.2,-1525.0,-746.07,-1193.3
1391.000000000,98.612,2269.0,2346.5,1814.9,338.20,3876.1,968.54,12.623,6199.2,2735.0,3367.1,2065.9,0.0000,-6574.7,-6877.5,-1227.3,-2033.8,-1867.7,-15431.,-102.48,-19117.,-6115.3,-3992.7,-2301.8,74.375,2649.6,2416.0,1886.7,373.69,4136.0,1686.6,0.0000,7310.7,4449.7,4252.8,3658.0,0.0000,-410.64,-125.89,-102.65,-49.583,-111.22,-587.69,0.0000,-1055.1,-1525.0,-746.05,-1193.2
1392.000000000,98.285,2259.5,2338.2,1808.6,336.82,3864.6,968.54,11.342,6189.6,2735.6,3366.8,2065.8,0.0000,-6574.9,-6876.1,-1227.2,-2033.2,-1868.2,-15430.,-102.44,-19116.,-6114.9,-3992.2,-2301.1,74.067,2638.6,2406.0,1878.3,372.14,4117.8,1686.6,0.0000,7299.7,4449.7,4252.8,3658.0,0.0000,-408.94,-125.35,-102.21,-49.378,-110.74,-587.69,0.0000,-1055.0,-1524.9,-746.04,-1193.1
1393.000000000,98.000,2249.9,2328.6,1802.3,335.50,3849.7,968.54,10.519,6179.7,2735.4,3366.8,2065.5,0.0000,-6574.6,-6874.5,-1227.0,-2032.7,-1868.6,-15429.,-102.40,-19116.,-6114.5,-3991.8,-2300.5,73.752,2627.4,2395.7,1869.7,370.54,4098.9,1686.6,0.0000,7288.3,4449.7,4252.8,3658.0,0.0000,-407.21,-124.80,-101.75,-49.168,-110.24,-587.69,0.0000,-1055.0,-1524.8,-746.03,-1193.0
1394.000000000,97.840,2240.1,2318.1,1794.6,334.08,3838.8,968.54,9.2882,6170.1,2735.0,3367.0,2065.3,0.0000,-6573.9,-6872.8,-1226.7,-2032.1,-1868.7,-15428.,-102.37,-19115.,-6114.1,-3991.4,-2299.9,73.433,2616.0,2385.4,1860.8,368.93,4079.4,1686.6,0.0000,7276.5,4449.7,4252.8,3658.0,0.0000,-405.44,-124.25,-101.28,-48.956,-109.73,-587.69,0.0000,-1054.9,-1524.8,-746.01,-1192.9
1395.000000000,97.695,2230.5,2307.5,1786.6,332.69,3822.5,968.54,9.2886,6165.6,2734.5,3366.8,2065.3,0.0000,-6572.7,-6870.9,-1226.4,-2031.5,-1868.7,-15426.,-102.33,-19115.,-6113.6,-3990.9,-2299.2,73.121,2604.9,2375.2,1851.9,367.34,4059.7,1686.6,0.0000,7264.6,4449.7,4252.8,3658.0,0.0000,-403.71,-123.69,-100.81,-48.747,-109.20,-587.69,0.0000,-1054.9,-1524.7,-746.00,-1192.8
1396.000000000,97.509,2221.2,2297.5,1778.3,331.29,3805.8,968.54,9.0556,6155.6,2734.2,3366.5,2065.5,0.0000,-6571.2,-6869.0,-1226.0,-2030.8,-1868.6,-15425.,-102.30,-19115.,-6113.2,-3990.5,-2298.6,72.808,2593.8,2365.1,1842.9,365.75,4039.8,1686.6,0.0000,7252.6,4449.7,4252.8,3658.0,0.0000,-401.97,-123.14,-100.34,-48.539,-108.66,-587.69,0.0000,-1054.8,-1524.7,-745.99,-1192.7
1397.000000000,97.193,2211.8,2287.7,1770.1,329.92,3794.0,968.54,7.9617,6148.2,2733.9,3366.8,2065.4,0.0000,-6569.3,-6866.9,-1225.5,-2030.2,-1868.3,-15424.,-102.26,-19114.,-6112.8,-3990.0,-2297.9,72.501,2582.8,2355.1,1833.8,364.19,4019.8,1686.6,0.0000,7240.5,4449.7,4252.8,3658.0,0.0000,-400.25,-122.59,-99.872,-48.334,-108.12,-587.69,0.0000,-1054.7,-1524.6,-745.97,-1192.6
1398.000000000,96.881,2202.6,2278.4,1761.9,328.56,3778.6,968.54,7.9622,6138.2,2733.7,3367.0,2065.3,0.0000,-6567.1,-6864.8,-1225.0,-2029.5,-1868.0,-15423.,-102.22,-19114.,-6112.3,-3989.6,-2297.3,72.202,2572.2,2345.4,1824.9,362.66,3999.9,1686.6,0.0000,7228.4,4449.7,4252.8,3658.0,0.0000,-398.57,-122.06,-99.409,-48.135,-107.57,-587.69,0.0000,-1054.7,-1524.5,-745.96,-1192.5
1399.000000000,96.602,2193.4,2269.3,1753.7,327.21,3762.8,968.55,7.9627,6127.9,2733.7,3367.0,2065.3,0.0000,-6564.6,-6862.7,-1224.4,-2028.8,-1867.5,-15421.,-102.19,-19113.,-6111.9,-3989.2,-2296.7,71.907,2561.6,2335.8,1815.9,361.15,3979.9,1686.6,0.0000,7216.3,4449.7,4252.8,3658.0,0.0000,-396.91,-121.53,-98.947,-47.938,-107.02,-587.69,0.0000,-1054.6,-1524.5,-745.95,-1192.4
1400.000000000,96.305,2184.5,2260.2,1745.3,325.88,3745.2,968.55,7.9632,6121.8,2733.3,3367.7,2065.3,0.0000,-6561.8,-6860.5,-1223.7,-2028.1,-1866.8,-15420.,-102.15,-19112.,-6111.4,-3988.7,-2296.0,71.615,2551.2,2326.3,1806.8,359.66,3959.7,1686.6,0.0000,7204.1,4449.7,4252.8,3658.0,0.0000,-395.26,-121.00,-98.484,-47.743,-106.46,-587.69,0.0000,-1054.5,-1524.4,-745.94,-1192.3
1401.000000000,95.765,2175.8,2250.6,1736.8,324.57,3727.5,968.51,7.9637,6114.4,2733.0,3367.9,2065.4,0.0000,-6558.8,-6858.2,-1223.0,-2027.3,-1866.1,-15419.,-102.12,-19111.,-6111.0,-3988.3,-2295.4,71.321,2540.8,2316.8,1797.7,358.15,3939.2,1686.6,0.0000,7191.7,4449.7,4252.8,3658.0,0.0000,-393.60,-120.47,-98.017,-47.547,-105.89,-587.69,0.0000,-1054.5,-1524.3,-745.92,-1192.2
1402.000000000,95.469,2166.9,2241.1,1728.4,323.25,3709.6,968.51,7.9642,6104.9,2732.9,3368.1,2065.5,0.0000,-6555.5,-6855.8,-1222.3,-2026.6,-1865.3,-15418.,-102.08,-19110.,-6110.5,-3987.9,-2294.8,71.018,2530.0,2306.9,1788.2,356.60,3918.1,1686.6,0.0000,7178.9,4449.7,4252.8,3658.0,0.0000,-391.88,-119.92,-97.533,-47.345,-105.30,-587.69,0.0000,-1054.4,-1524.3,-745.91,-1192.1
1403.000000000,95.182,2157.8,2231.8,1719.8,321.94,3694.4,968.51,7.9647,6093.9,2732.8,3368.5,2065.5,0.0000,-6552.0,-6853.3,-1221.5,-2025.8,-1864.3,-15416.,-102.05,-19109.,-6110.1,-3987.4,-2294.1,70.724,2519.5,2297.4,1778.9,355.09,3897.2,1686.6,0.0000,7166.3,4449.7,4252.8,3658.0,0.0000,-390.22,-119.38,-97.060,-47.150,-104.71,-587.69,0.0000,-1054.3,-1524.2,-745.90,-1192.0
1404.000000000,94.850,2153.5,2226.9,1712.9,321.44,3678.0,968.51,7.4052,6083.3,2732.7,3368.6,2065.6,0.0000,-6548.6,-6851.0,-1220.7,-2025.1,-1863.3,-15415.,-102.01,-19108.,-6109.6,-3987.0,-2293.5,79.304,2569.4,2337.4,1811.2,372.45,3935.4,1686.6,9.9293,7199.9,4461.4,4265.9,3670.0,0.0000,-393.73,-120.84,-97.777,-47.662,-105.39,-587.69,-0.45336,-1054.6,-1524.2,-745.95,-1192.1
1405.000000000,95.198,2157.9,2229.7,1709.4,322.12,3666.3,968.51,6.6378,6073.8,2732.6,3368.5,2065.5,0.0000,-6546.0,-6849.1,-1219.9,-2024.4,-1862.4,-15414.,-101.98,-19107.,-6109.2,-3986.6,-2292.9,71.438,2544.9,2320.6,1785.2,358.48,3905.4,1686.6,0.0000,7171.1,4449.7,4252.8,3658.0,0.0000,-394.07,-120.52,-97.629,-47.625,-104.90,-587.69,0.0000,-1054.3,-1524.1,-745.87,-1191.8
1406.000000000,95.214,2159.2,2231.7,1706.5,322.16,3655.8,968.51,6.6545,6065.2,2732.3,3368.6,2065.6,0.0000,-6543.7,-6847.5,-1219.2,-2023.8,-1861.5,-15413.,-101.94,-19106.,-6108.7,-3986.1,-2292.3,71.291,2539.7,2315.8,1777.3,357.67,3886.5,1686.6,0.0000,7159.7,4449.7,4252.8,3658.0,0.0000,-393.22,-120.25,-97.278,-47.527,-104.36,-587.69,0.0000,-1054.2,-1524.0,-745.86,-1191.7
1407.000000000,95.257,2156.9,2229.0,1702.6,322.33,3642.8,968.51,6.6668,6056.1,2732.3,3368.3,2065.5,0.0000,-6541.4,-6845.8,-1218.4,-2023.1,-1860.6,-15411.,-101.91,-19105.,-6108.3,-3985.7,-2291.6,71.182,2535.8,2312.3,1770.9,357.06,3871.1,1686.6,0.0000,7150.3,4449.7,4252.8,3658.0,0.0000,-392.58,-120.04,-96.998,-47.455,-103.91,-587.69,0.0000,-1054.2,-1524.0,-745.85,-1191.6
1408.000000000,95.239,2154.6,2225.0,1698.7,321.86,3628.5,968.51,5.8735,6046.5,2732.2,3367.8,2065.5,0.0000,-6539.0,-6844.1,-1217.6,-2022.4,-1859.5,-15410.,-101.87,-19104.,-6107.8,-3985.3,-2291.0,70.951,2527.6,2304.7,1762.1,355.84,3850.8,1686.6,0.0000,7138.0,4449.7,4252.8,3658.0,0.0000,-391.26,-119.62,-96.573,-47.300,-103.33,-587.69,0.0000,-1054.1,-1523.9,-745.84,-1191.5
1409.000000000,94.953,2150.7,2219.6,1694.4,321.03,3612.7,968.51,5.3562,6037.6,2732.1,3367.5,2065.7,0.0000,-6536.3,-6842.3,-1216.9,-2021.8,-1858.3,-15409.,-101.84,-19102.,-6107.3,-3984.9,-2290.4,70.727,2519.6,2297.5,1753.5,354.67,3831.2,1686.6,0.0000,7126.2,4449.7,4252.8,3658.0,0.0000,-389.99,-119.21,-96.162,-47.151,-102.77,-587.69,0.0000,-1054.0,-1523.9,-745.82,-1191.4
1410.000000000,94.750,2151.7,2220.5,1688.1,321.35,3599.1,968.51,5.3568,6030.8,2732.1,3367.5,2065.6,0.0000,-6534.1,-6840.8,-1216.1,-2021.1,-1857.0,-15407.,-101.80,-19101.,-6106.9,-3984.4,-2289.8,107.33,2719.5,2440.7,1806.7,386.53,3888.5,1686.6,36.889,7176.5,4469.6,4274.7,3678.4,0.0000,-396.78,-123.43,-97.345,-48.106,-103.69,-587.69,-1.6843,-1054.5,-1523.8,-745.92,-1191.6
1411.000000000,95.296,2165.6,2232.7,1684.5,323.41,3595.3,968.51,5.3575,6026.1,2732.0,3367.4,2065.8,0.0000,-6533.0,-6840.0,-1215.4,-2020.6,-1855.8,-15406.,-101.77,-19100.,-6106.4,-3984.0,-2289.2,72.270,2574.6,2347.6,1767.4,362.18,3848.7,1686.6,0.0000,7136.5,4449.7,4252.8,3658.0,0.0000,-398.45,-121.78,-97.400,-48.181,-103.18,-587.69,0.0000,-1054.0,-1523.7,-745.80,-1191.2
1412.000000000,95.551,2175.2,2242.2,1683.7,324.38,3591.5,968.51,5.3582,6020.9,2732.0,3367.8,2065.7,0.0000,-6532.6,-6839.6,-1214.7,-2020.1,-1854.7,-15405.,-101.73,-19099.,-6106.0,-3983.6,-2288.6,72.251,2573.9,2347.0,1759.8,361.79,3830.4,1686.6,0.0000,7125.3,4449.7,4252.8,3658.0,0.0000,-398.32,-121.74,-97.142,-48.167,-102.65,-587.69,0.0000,-1053.9,-1523.7,-745.79,-1191.1
1413.000000000,95.833,2178.0,2245.3,1682.2,325.39,3581.1,968.52,5.3612,6013.8,2731.9,3368.2,2065.7,0.0000,-6532.3,-6839.2,-1214.0,-2019.6,-1853.5,-15403.,-101.70,-19097.,-6105.5,-3983.1,-2288.1,72.139,2569.9,2343.3,1752.1,361.13,3811.6,1686.6,0.0000,7113.9,4449.7,4252.8,3658.0,0.0000,-397.69,-121.54,-96.816,-48.093,-102.11,-587.69,0.0000,-1053.9,-1523.6,-745.77,-1191.0
1414.000000000,95.952,2176.9,2245.4,1678.8,325.26,3568.0,968.52,5.3692,6005.5,2731.8,3368.4,2065.7,0.0000,-6531.7,-6838.6,-1213.2,-2019.1,-1852.2,-15402.,-101.66,-19096.,-6105.1,-3982.7,-2287.5,71.979,2564.2,2338.1,1744.1,360.25,3792.6,1686.6,0.0000,7102.4,4449.7,4252.8,3658.0,0.0000,-396.79,-121.26,-96.455,-47.986,-101.56,-587.69,0.0000,-1053.8,-1523.5,-745.76,-1190.9
1415.000000000,95.701,2174.2,2242.6,1673.4,324.54,3553.1,968.52,5.3698,5997.3,2731.7,3368.5,2065.6,0.0000,-6530.8,-6837.9,-1212.4,-2018.5,-1850.8,-15400.,-101.63,-19094.,-6104.6,-3982.3,-2287.0,71.792,2557.5,2332.0,1735.9,359.25,3773.4,1686.6,0.0000,7090.8,4449.7,4252.8,3658.0,0.0000,-395.74,-120.94,-96.074,-47.861,-101.00,-587.69,0.0000,-1053.7,-1523.5,-745.75,-1190.8
1416.000000000,95.547,2169.9,2238.6,1666.9,323.64,3538.4,968.52,5.2341,5992.0,2731.7,3368.3,2065.7,0.0000,-6529.6,-6837.1,-1211.6,-2017.9,-1849.2,-15399.,-101.59,-19093.,-6104.2,-3981.8,-2286.4,71.585,2550.2,2325.3,1727.6,358.16,3754.1,1686.6,0.0000,7079.1,4449.7,4252.8,3658.0,0.0000,-394.58,-120.58,-95.677,-47.723,-100.44,-587.69,0.0000,-1053.7,-1523.4,-745.74,-1190.7
1417.000000000,95.360,2165.4,2234.8,1659.4,322.77,3526.6,968.52,4.0431,5988.6,2731.7,3368.2,2065.7,0.0000,-6528.1,-6836.1,-1210.7,-2017.3,-1847.6,-15398.,-101.56,-19092.,-6103.7,-3981.4,-2285.9,71.365,2542.3,2318.2,1719.1,357.01,3734.7,1686.6,0.0000,7067.3,4449.7,4252.8,3658.0,0.0000,-393.35,-120.19,-95.270,-47.577,-99.868,-587.69,0.0000,-1053.6,-1523.4,-745.72,-1190.6
1418.000000000,95.152,2160.4,2230.0,1652.9,321.79,3514.6,968.52,4.0439,5981.3,2731.7,3368.1,2065.9,0.0000,-6526.5,-6835.0,-1209.7,-2016.7,-1845.9,-15396.,-101.52,-19090.,-6103.3,-3981.0,-2285.4,71.137,2534.2,2310.8,1710.6,355.82,3715.2,1686.6,0.0000,7055.5,4449.7,4252.8,3658.0,0.0000,-392.07,-119.79,-94.856,-47.424,-99.293,-587.69,0.0000,-1053.5,-1523.3,-745.71,-1190.5
1419.000000000,94.932,2154.7,2223.8,1648.4,320.80,3499.1,968.52,4.0447,5972.4,2731.7,3368.0,2066.0,0.0000,-6524.5,-6833.8,-1208.6,-2016.0,-1844.1,-15395.,-101.49,-19089.,-6102.8,-3980.6,-2284.9,70.943,2527.3,2304.5,1702.9,354.79,3697.3,1686.6,0.0000,7044.6,4449.7,4252.8,3658.0,0.0000,-390.97,-119.44,-94.486,-47.295,-98.761,-587.69,0.0000,-1053.4,-1523.2,-745.70,-1190.4
1420.000000000,94.724,2150.1,2217.9,1641.5,319.83,3482.3,968.52,4.0454,5962.8,2731.7,3368.0,2066.1,0.0000,-6522.4,-6832.5,-1207.5,-2015.3,-1842.3,-15394.,-101.45,-19087.,-6102.3,-3980.1,-2284.3,70.754,2520.6,2298.3,1695.4,353.80,3679.8,1686.6,0.0000,7034.0,4449.7,4252.8,3658.0,0.0000,-389.90,-119.10,-94.124,-47.169,-98.238,-587.69,0.0000,-1053.4,-1523.2,-745.69,-1190.3
1421.000000000,94.520,2145.3,2212.9,1634.1,318.87,3465.6,968.52,4.0462,5952.5,2731.7,3367.9,2066.0,0.0000,-6520.0,-6831.1,-1206.4,-2014.6,-1840.4,-15392.,-101.41,-19086.,-6101.9,-3979.7,-2283.8,70.555,2513.5,2291.9,1687.6,352.75,3661.9,1686.6,0.0000,7023.2,4449.7,4252.8,3658.0,0.0000,-388.77,-118.74,-93.750,-47.036,-97.704,-587.69,0.0000,-1053.3,-1523.1,-745.67,-1190.2
1422.000000000,94.318,2139.5,2206.8,1626.8,317.99,3449.4,968.52,4.0510,5942.2,2731.6,3367.7,2066.0,0.0000,-6517.3,-6829.7,-1205.2,-2013.9,-1838.4,-15391.,-101.38,-19084.,-6101.4,-3979.3,-2283.3,70.341,2505.9,2284.9,1679.6,351.63,3643.6,1686.6,0.0000,7012.1,4449.7,4252.8,3658.0,0.0000,-387.55,-118.36,-93.361,-46.894,-97.155,-587.69,0.0000,-1053.2,-1523.0,-745.66,-1190.1
1423.000000000,94.111,2133.9,2200.7,1619.4,317.04,3434.1,968.52,4.0616,5932.4,2731.5,3367.5,2066.0,0.0000,-6514.5,-6828.2,-1204.0,-2013.2,-1836.4,-15389.,-101.34,-19083.,-6101.0,-3978.8,-2282.8,70.118,2497.9,2277.7,1671.5,350.47,3624.9,1686.6,0.0000,7000.8,4449.7,4252.8,3658.0,0.0000,-386.29,-117.96,-92.960,-46.745,-96.594,-587.69,0.0000,-1053.2,-1523.0,-745.65,-1190.0
1424.000000000,93.896,2127.8,2194.9,1612.2,316.06,3420.1,968.53,4.0624,5922.3,2731.6,3367.4,2066.1,0.0000,-6511.5,-6826.7,-1202.8,-2012.5,-1834.4,-15388.,-101.31,-19081.,-6100.5,-3978.4,-2282.2,69.907,2490.4,2270.8,1663.6,349.37,3606.8,1686.6,0.0000,6989.8,4449.7,4252.8,3658.0,0.0000,-385.08,-117.58,-92.575,-46.605,-96.048,-587.69,0.0000,-1053.1,-1522.9,-745.64,-1189.9
1425.000000000,93.829,2121.9,2188.8,1604.9,315.08,3406.5,968.53,4.0632,5912.4,2731.6,3367.3,2066.2,0.0000,-6508.4,-6825.0,-1201.6,-2011.7,-1832.3,-15386.,-101.27,-19080.,-6100.1,-3978.0,-2281.7,69.691,2482.7,2263.8,1655.6,348.24,3588.5,1686.6,0.0000,6978.8,4449.7,4252.8,3658.0,0.0000,-383.85,-117.18,-92.184,-46.461,-95.495,-587.69,0.0000,-1053.0,-1522.9,-745.63,-1189.8
1426.000000000,93.650,2116.3,2182.5,1597.6,314.14,3390.3,968.53,4.0639,5902.7,2731.5,3367.3,2066.1,0.0000,-6505.1,-6823.2,-1200.3,-2011.0,-1830.1,-15385.,-101.24,-19078.,-6099.6,-3977.5,-2281.2,69.537,2477.2,2258.8,1650.9,348.18,3578.0,1686.6,0.0000,6972.4,4449.7,4252.8,3658.0,0.0000,-382.95,-116.89,-91.935,-46.362,-95.154,-587.69,0.0000,-1052.9,-1522.8,-745.61,-1189.7
1427.000000000,93.465,2110.8,2177.1,1590.6,313.27,3376.7,968.53,4.0646,5893.1,2731.5,3367.1,2066.1,0.0000,-6501.7,-6821.5,-1199.0,-2010.2,-1827.9,-15384.,-101.20,-19076.,-6099.2,-3977.1,-2280.7,69.325,2469.7,2251.9,1643.0,346.34,3559.9,1686.6,0.0000,6961.4,4449.7,4252.8,3658.0,0.0000,-381.74,-116.51,-91.549,-46.216,-94.604,-587.69,0.0000,-1052.9,-1522.7,-745.60,-1189.6
1428.000000000,93.257,2104.8,2171.2,1584.2,312.36,3363.0,968.53,4.0654,5883.7,2731.9,3367.0,2066.2,0.0000,-6498.2,-6819.6,-1197.6,-2009.4,-1825.8,-15382.,-101.17,-19075.,-6098.8,-3976.7,-2280.1,69.103,2461.8,2244.7,1634.9,345.19,3541.4,1686.6,0.0000,6950.3,4449.7,4252.8,3658.0,0.0000,-380.47,-116.10,-91.152,-46.069,-94.043,-587.69,0.0000,-1052.8,-1522.7,-745.59,-1189.5
1429.000000000,93.048,2098.5,2164.9,1577.6,311.49,3347.0,968.52,4.0661,5873.9,2732.3,3367.0,2066.2,0.0000,-6494.6,-6817.7,-1196.3,-2008.6,-1823.5,-15381.,-101.13,-19073.,-6098.3,-3976.2,-2279.6,68.898,2454.4,2238.0,1627.2,344.11,3523.6,1686.6,0.0000,6939.5,4449.7,4252.8,3658.0,0.0000,-379.28,-115.72,-90.774,-45.932,-93.504,-587.69,0.0000,-1052.7,-1522.6,-745.58,-1189.4
1430.000000000,92.574,2092.5,2159.1,1570.8,310.53,3331.4,968.50,4.0668,5864.0,2732.3,3367.3,2066.3,0.0000,-6490.8,-6815.8,-1194.9,-2007.8,-1821.2,-15379.,-101.10,-19071.,-6097.9,-3975.8,-2279.1,68.695,2447.2,2231.5,1619.5,343.05,3506.0,1686.6,0.0000,6928.8,4449.7,4252.8,3658.0,0.0000,-378.11,-115.35,-90.400,-45.797,-92.979,-587.69,0.0000,-1052.6,-1522.6,-745.56,-1189.3
1431.000000000,92.364,2086.5,2153.1,1563.8,309.60,3315.4,968.47,4.0676,5854.5,2732.2,3367.2,2066.2,0.0000,-6486.9,-6813.8,-1193.5,-2007.0,-1818.8,-15378.,-101.06,-19070.,-6097.4,-3975.4,-2278.6,68.512,2440.7,2225.5,1612.2,342.08,3489.1,1686.6,0.0000,6918.6,4449.7,4252.8,3658.0,0.0000,-377.05,-115.00,-90.049,-45.674,-92.474,-587.69,0.0000,-1052.6,-1522.5,-745.55,-1189.2
1432.000000000,92.097,2080.8,2147.8,1556.7,308.70,3299.4,968.47,4.0683,5845.2,2732.3,3367.2,2066.3,0.0000,-6483.0,-6811.8,-1192.1,-2006.2,-1816.4,-15376.,-101.03,-19068.,-6097.0,-3974.9,-2278.1,68.324,2434.0,2219.4,1604.9,341.10,3472.1,1686.6,0.0000,6908.3,4449.7,4252.8,3658.0,0.0000,-375.96,-114.65,-89.693,-45.549,-91.965,-587.69,0.0000,-1052.5,-1522.4,-745.54,-1189.1
1433.000000000,91.698,2077.5,2144.8,1549.7,308.21,3284.8,968.47,4.0690,5836.1,2732.3,3367.2,2066.3,0.0000,-6479.2,-6809.8,-1190.7,-2005.4,-1813.9,-15375.,-100.99,-19066.,-6096.5,-3974.5,-2277.5,78.232,2453.4,2241.2,1605.8,345.68,3468.5,1686.6,1.6541,6906.6,4450.6,4253.5,3658.7,0.0000,-377.54,-115.37,-89.827,-45.767,-91.805,-587.69,-0.75525E-01,-1052.5,-1522.4,-745.53,-1189.0
1434.000000000,91.831,2082.4,2148.3,1544.0,309.06,3272.6,968.47,4.0697,5827.5,2732.3,3367.1,2066.4,0.0000,-6476.0,-6808.2,-1189.3,-2004.7,-1811.5,-15373.,-100.96,-19065.,-6096.1,-3974.1,-2277.0,118.67,2545.8,2316.6,1625.8,361.68,3489.6,1686.6,23.905,6923.3,4457.1,4260.2,3665.2,0.0000,-382.00,-117.74,-90.522,-46.375,-92.147,-587.69,-1.0915,-1052.6,-1522.3,-745.55,-1189.1
1435.000000000,92.367,2119.6,2181.6,1542.5,315.21,3267.7,968.47,4.0705,5820.2,2732.3,3367.0,2066.4,0.0000,-6475.9,-6808.5,-1188.4,-2004.3,-1809.3,-15372.,-100.93,-19063.,-6095.7,-3973.6,-2276.5,832.51,3837.2,3219.7,1718.2,416.00,3624.7,1686.6,576.46,7013.2,4477.5,4280.5,3685.4,0.0000,-413.46,-142.34,-95.555,-50.147,-95.209,-587.69,-26.321,-1053.1,-1522.2,-745.64,-1189.3
1436.000000000,95.417,2197.1,2249.6,1550.9,326.81,3276.0,968.47,4.0712,5816.9,2732.1,3367.0,2066.5,0.0000,-6481.0,-6811.8,-1187.7,-2004.5,-1807.5,-15370.,-100.90,-19061.,-6095.3,-3973.2,-2276.0,249.77,2834.6,2630.0,1807.4,452.95,3644.8,1686.8,0.0000,7050.8,4491.5,4289.1,3691.1,0.0000,-419.71,-131.23,-96.431,-51.292,-95.124,-587.69,0.0000,-1053.6,-1522.2,-745.67,-1189.3
1437.000000000,97.067,2249.3,2305.3,1567.3,333.86,3286.4,968.43,4.0719,5815.3,2732.2,3367.0,2066.7,0.0000,-6488.6,-6816.7,-1187.3,-2004.9,-1806.1,-15369.,-100.87,-19060.,-6094.8,-3972.8,-2275.5,77.272,2752.8,2510.1,1749.8,406.42,3610.4,1686.6,0.0000,7020.8,4482.2,4278.2,3681.3,0.0000,-425.20,-129.75,-96.923,-51.656,-94.618,-587.69,0.0000,-1053.3,-1522.1,-745.60,-1189.0
1438.000000000,99.175,2281.5,2336.8,1577.8,341.71,3288.7,968.42,4.0727,5812.6,2732.2,3367.1,2067.0,0.0000,-6497.2,-6821.5,-1186.9,-2005.3,-1804.7,-15367.,-100.84,-19058.,-6094.4,-3972.3,-2275.0,77.460,2759.5,2516.2,1726.2,403.55,3589.0,1686.6,0.0000,6999.1,4476.2,4274.0,3677.6,0.0000,-426.32,-130.14,-96.849,-51.759,-94.151,-587.69,0.0000,-1053.0,-1522.1,-745.57,-1188.9
1439.000000000,100.28,2296.8,2356.4,1583.6,343.81,3285.0,968.42,4.0525,5808.7,2732.3,3367.1,2067.2,0.0000,-6505.5,-6825.8,-1186.5,-2005.6,-1803.1,-15366.,-100.80,-19056.,-6094.0,-3971.9,-2274.5,77.464,2759.6,2516.3,1708.6,399.29,3568.4,1686.6,0.0000,6980.0,4468.8,4269.0,3672.9,0.0000,-426.44,-130.22,-96.663,-51.736,-93.705,-587.69,0.0000,-1052.8,-1522.0,-745.54,-1188.7
1440.000000000,100.67,2304.3,2364.4,1584.5,344.52,3280.5,968.43,3.5313,5808.1,2732.3,3367.3,2067.2,0.0000,-6512.9,-6829.6,-1186.2,-2005.7,-1801.3,-15364.,-100.77,-19055.,-6093.6,-3971.4,-2273.9,77.369,2756.2,2513.2,1689.8,394.03,3546.0,1686.6,0.0000,6961.3,4462.4,4263.1,3667.4,0.0000,-426.02,-130.14,-96.406,-51.643,-93.242,-587.69,0.0000,-1052.6,-1521.9,-745.49,-1188.5
1441.000000000,100.71,2307.3,2370.4,1583.3,344.22,3275.1,968.43,3.5319,5809.8,2732.3,3367.5,2067.2,0.0000,-6519.6,-6832.9,-1185.7,-2005.7,-1799.3,-15363.,-100.73,-19053.,-6093.2,-3971.0,-2273.4,77.209,2750.5,2508.0,1675.7,389.40,3526.4,1686.6,0.0000,6945.5,4457.7,4259.9,3664.4,0.0000,-425.23,-129.94,-96.099,-51.513,-92.778,-587.69,0.0000,-1052.4,-1521.9,-745.47,-1188.4
1442.000000000,100.61,2307.8,2374.6,1578.7,343.59,3274.4,968.43,3.5326,5816.6,2732.4,3367.4,2067.3,0.0000,-6525.7,-6835.6,-1185.0,-2005.7,-1797.2,-15361.,-100.70,-19051.,-6092.7,-3970.6,-2272.9,77.002,2743.1,2501.3,1662.8,385.52,3506.8,1686.6,0.0000,6931.4,4454.3,4256.9,3661.7,0.0000,-424.18,-129.65,-95.749,-51.357,-92.296,-587.69,0.0000,-1052.3,-1521.8,-745.44,-1188.3
1443.000000000,100.59,2308.5,2375.1,1574.4,342.78,3275.3,968.43,3.5332,5819.2,2732.3,3367.5,2067.4,0.0000,-6531.2,-6837.9,-1184.3,-2005.5,-1795.1,-15360.,-100.67,-19050.,-6092.3,-3970.1,-2272.4,76.813,2736.4,2495.2,1652.4,382.65,3490.3,1686.6,0.0000,6919.5,4452.1,4254.9,3659.9,0.0000,-423.23,-129.38,-95.438,-51.220,-91.872,-587.69,0.0000,-1052.2,-1521.8,-745.42,-1188.1
1444.000000000,100.45,2305.4,2371.4,1571.9,341.87,3269.7,968.43,3.5339,5816.7,2732.3,3367.4,2067.5,0.0000,-6535.9,-6839.8,-1183.4,-2005.3,-1792.9,-15358.,-100.63,-19048.,-6091.9,-3969.7,-2271.9,76.568,2727.7,2487.2,1644.2,380.58,3473.4,1686.6,0.0000,6909.1,4451.4,4254.2,3659.2,0.0000,-421.95,-129.01,-95.059,-51.052,-91.393,-587.69,0.0000,-1052.1,-1521.7,-745.40,-1188.0
1445.000000000,100.22,2303.6,2366.5,1568.8,340.86,3258.4,968.43,3.5345,5810.9,2732.3,3367.4,2067.6,0.0000,-6539.8,-6841.4,-1182.5,-2005.1,-1790.6,-15357.,-100.60,-19047.,-6091.5,-3969.3,-2271.4,76.323,2719.0,2479.2,1634.9,378.70,3456.5,1686.6,0.0000,6897.8,4450.4,4253.4,3658.5,0.0000,-420.66,-128.64,-94.683,-50.884,-90.920,-587.69,0.0000,-1052.0,-1521.6,-745.39,-1187.9
1446.000000000,99.989,2300.5,2363.2,1563.6,339.83,3247.3,968.43,3.5352,5803.7,2732.3,3367.4,2067.7,0.0000,-6542.8,-6842.9,-1181.5,-2004.8,-1788.4,-15355.,-100.56,-19045.,-6091.1,-3968.8,-2270.9,76.094,2710.8,2471.8,1627.2,377.26,3441.3,1686.6,0.0000,6888.2,4450.0,4253.0,3658.2,0.0000,-419.46,-128.29,-94.332,-50.730,-90.478,-587.69,0.0000,-1051.9,-1521.6,-745.37,-1187.8
1447.000000000,99.697,2295.2,2359.0,1557.4,338.75,3234.1,968.38,3.5358,5795.6,2732.3,3367.4,2067.7,0.0000,-6545.1,-6844.1,-1180.5,-2004.5,-1786.0,-15354.,-100.53,-19043.,-6090.7,-3968.4,-2270.3,75.830,2701.4,2463.2,1619.5,375.85,3425.0,1686.6,0.0000,6878.2,4449.8,4252.9,3658.1,0.0000,-418.05,-127.87,-93.940,-50.554,-90.000,-587.69,0.0000,-1051.9,-1521.5,-745.36,-1187.7
1448.000000000,99.331,2290.7,2354.1,1551.1,337.66,3222.2,968.35,3.5364,5788.0,2732.4,3367.3,2067.8,0.0000,-6547.1,-6845.1,-1179.4,-2004.2,-1783.7,-15352.,-100.49,-19042.,-6090.2,-3967.9,-2269.8,75.587,2692.8,2455.3,1612.4,374.57,3409.7,1686.6,0.0000,6868.9,4449.7,4252.8,3658.0,0.0000,-416.76,-127.48,-93.573,-50.391,-89.545,-587.69,0.0000,-1051.8,-1521.5,-745.35,-1187.6
1449.000000000,99.137,2284.5,2350.7,1544.7,336.67,3210.7,968.35,3.5371,5781.2,2732.4,3367.4,2067.9,0.0000,-6548.8,-6845.8,-1178.3,-2003.8,-1781.3,-15351.,-100.46,-19040.,-6089.8,-3967.5,-2269.3,75.398,2686.0,2449.2,1606.5,373.59,3396.5,1686.6,0.0000,6860.8,4449.7,4252.8,3658.0,0.0000,-415.75,-127.18,-93.267,-50.265,-89.143,-587.69,0.0000,-1051.7,-1521.4,-745.33,-1187.6
1450.000000000,98.491,2280.4,2345.1,1539.0,335.70,3198.8,968.35,3.5389,5773.1,2732.4,3367.3,2068.0,0.0000,-6550.1,-6846.4,-1177.2,-2003.4,-1778.9,-15349.,-100.42,-19038.,-6089.4,-3967.1,-2268.8,75.192,2678.7,2442.5,1600.3,372.54,3382.7,1686.6,0.0000,6852.5,4449.7,4252.8,3658.0,0.0000,-414.65,-126.85,-92.944,-50.128,-88.727,-587.69,0.0000,-1051.6,-1521.3,-745.32,-1187.5
1451.000000000,98.527,2275.0,2338.7,1533.3,334.77,3186.3,968.36,3.5442,5764.8,2732.4,3367.2,2068.0,0.0000,-6551.0,-6846.7,-1176.0,-2003.0,-1776.5,-15347.,-100.39,-19037.,-6089.0,-3966.6,-2268.3,74.955,2670.2,2434.8,1593.6,371.34,3368.0,1686.6,0.0000,6843.6,4449.7,4252.8,3658.0,0.0000,-413.36,-126.46,-92.586,-49.970,-88.283,-587.69,0.0000,-1051.6,-1521.3,-745.31,-1187.4
1452.000000000,98.321,2268.7,2332.0,1527.4,333.80,3172.9,968.32,3.5448,5757.5,2732.4,3367.3,2068.1,0.0000,-6551.5,-6846.8,-1174.8,-2002.6,-1774.1,-15346.,-100.36,-19035.,-6088.6,-3966.2,-2267.8,74.746,2662.8,2428.0,1587.6,370.28,3354.8,1686.6,0.0000,6835.7,4449.7,4252.8,3658.0,0.0000,-412.24,-126.12,-92.268,-49.831,-87.882,-587.69,0.0000,-1051.5,-1521.2,-745.30,-1187.3
1453.000000000,98.116,2262.5,2325.3,1522.3,332.72,3159.8,968.32,3.4835,5749.8,2732.5,3367.3,2068.2,0.0000,-6551.7,-6846.7,-1173.6,-2002.1,-1771.6,-15344.,-100.32,-19033.,-6088.2,-3965.7,-2267.3,74.497,2653.9,2419.9,1580.7,369.02,3339.7,1686.6,0.0000,6826.5,4449.7,4252.8,3658.0,0.0000,-410.88,-125.70,-91.897,-49.665,-87.426,-587.69,0.0000,-1051.4,-1521.2,-745.29,-1187.2
1454.000000000,97.708,2256.7,2318.5,1516.7,331.74,3148.1,968.32,3.0316,5742.2,2732.5,3367.3,2068.3,0.0000,-6551.4,-6846.4,-1172.3,-2001.6,-1769.2,-15343.,-100.29,-19031.,-6087.8,-3965.3,-2266.8,74.339,2648.3,2414.8,1575.5,368.20,3327.9,1686.6,0.0000,6819.4,4449.7,4252.8,3658.0,0.0000,-410.01,-125.43,-91.631,-49.559,-87.061,-587.69,0.0000,-1051.4,-1521.1,-745.27,-1187.1
1455.000000000,97.150,2251.4,2311.8,1511.7,330.84,3137.5,968.32,3.0322,5734.3,2732.7,3367.2,2068.4,0.0000,-6550.9,-6845.9,-1171.0,-2001.1,-1766.7,-15341.,-100.25,-19030.,-6087.3,-3964.8,-2266.2,74.069,2638.7,2406.0,1568.2,366.84,3312.1,1686.6,0.0000,6809.8,4449.7,4252.8,3658.0,0.0000,-408.53,-124.97,-91.237,-49.380,-86.586,-587.69,0.0000,-1051.3,-1521.0,-745.26,-1187.0
1456.000000000,96.886,2244.2,2305.8,1506.5,329.74,3125.2,968.32,3.0328,5726.9,2732.7,3367.3,2068.4,0.0000,-6550.0,-6845.3,-1169.7,-2000.6,-1764.2,-15340.,-100.22,-19028.,-6086.9,-3964.4,-2265.7,73.794,2628.9,2397.1,1560.9,365.45,3296.0,1686.6,0.0000,6800.1,4449.7,4252.8,3658.0,0.0000,-407.01,-124.50,-90.836,-49.196,-86.105,-587.69,0.0000,-1051.2,-1521.0,-745.25,-1186.9
1457.000000000,96.588,2236.6,2301.6,1500.3,328.63,3112.6,968.32,3.0334,5720.2,2733.1,3367.4,2068.5,0.0000,-6548.9,-6844.4,-1168.4,-2000.0,-1761.6,-15338.,-100.18,-19026.,-6086.5,-3964.0,-2265.2,73.526,2619.3,2388.4,1553.6,364.09,3280.2,1686.6,0.0000,6790.5,4449.7,4252.8,3658.0,0.0000,-405.52,-124.03,-90.444,-49.017,-85.631,-587.69,0.0000,-1051.1,-1520.9,-745.24,-1186.8
1458.000000000,96.353,2229.9,2296.1,1494.0,327.40,3099.3,968.28,3.0340,5713.8,2733.5,3367.4,2068.5,0.0000,-6547.7,-6843.4,-1167.0,-1999.4,-1759.0,-15337.,-100.15,-19024.,-6086.1,-3963.5,-2264.7,73.259,2609.8,2379.7,1546.4,362.74,3264.4,1686.6,0.0000,6781.0,4449.7,4252.8,3658.0,0.0000,-404.04,-123.56,-90.053,-48.839,-85.157,-587.69,0.0000,-1051.1,-1520.9,-745.22,-1186.7
1459.000000000,96.116,2222.4,2288.8,1487.7,326.22,3088.8,968.28,3.0346,5706.0,2733.5,3367.4,2068.6,0.0000,-6546.1,-6842.1,-1165.6,-1998.8,-1756.3,-15335.,-100.12,-19023.,-6085.7,-3963.1,-2264.2,72.992,2600.3,2371.0,1539.2,361.39,3248.7,1686.6,0.0000,6771.4,4449.7,4252.8,3658.0,0.0000,-402.55,-123.09,-89.661,-48.661,-84.682,-587.69,0.0000,-1051.0,-1520.8,-745.21,-1186.6
1460.000000000,95.590,2215.3,2282.5,1482.2,325.10,3075.7,968.28,3.0351,5698.5,2733.6,3367.3,2068.6,0.0000,-6544.4,-6840.8,-1164.2,-1998.2,-1753.6,-15333.,-100.08,-19021.,-6085.3,-3962.6,-2263.7,72.788,2593.0,2364.4,1533.0,360.35,3235.0,1686.6,0.0000,6763.2,4449.7,4252.8,3658.0,0.0000,-401.40,-122.73,-89.340,-48.525,-84.264,-587.69,0.0000,-1050.9,-1520.7,-745.20,-1186.5
1461.000000000,95.382,2208.3,2278.5,1476.1,324.08,3062.7,968.28,3.0929,5690.5,2733.8,3367.4,2068.7,0.0000,-6542.6,-6839.4,-1162.7,-1997.5,-1750.9,-15332.,-100.05,-19019.,-6084.9,-3962.2,-2263.2,72.564,2585.0,2357.1,1526.6,359.22,3220.8,1686.6,0.0000,6754.6,4449.7,4252.8,3658.0,0.0000,-400.14,-122.33,-88.997,-48.376,-83.831,-587.69,0.0000,-1050.9,-1520.7,-745.19,-1186.4
1462.000000000,95.151,2201.6,2272.6,1469.9,323.06,3049.5,968.24,5.0082,5682.2,2733.8,3367.4,2068.7,0.0000,-6540.6,-6837.9,-1161.2,-1996.9,-1748.2,-15330.,-100.01,-19017.,-6084.5,-3961.8,-2262.7,72.321,2576.4,2349.2,1519.8,357.98,3206.0,1686.6,0.0000,6745.6,4449.7,4252.8,3658.0,0.0000,-398.77,-121.89,-88.634,-48.214,-83.380,-587.69,0.0000,-1050.8,-1520.6,-745.18,-1186.3
1463.000000000,94.916,2194.7,2265.8,1463.7,322.05,3036.9,968.25,5.0132,5673.9,2733.8,3367.4,2068.8,0.0000,-6538.3,-6836.3,-1159.7,-1996.2,-1745.4,-15329.,-99.978,-19015.,-6084.1,-3961.3,-2262.2,72.127,2569.5,2342.9,1513.4,356.98,3191.6,1686.6,0.0000,6736.9,4449.7,4252.8,3658.0,0.0000,-397.67,-121.54,-88.309,-48.084,-82.942,-587.69,0.0000,-1050.7,-1520.6,-745.16,-1186.2
1464.000000000,94.705,2188.4,2258.8,1457.5,321.12,3023.6,968.25,5.0179,5665.5,2733.8,3367.3,2068.9,0.0000,-6535.9,-6834.6,-1158.2,-1995.5,-1742.6,-15327.,-99.945,-19013.,-6083.7,-3960.9,-2261.7,71.890,2561.0,2335.2,1506.8,355.78,3177.0,1686.6,0.0000,6728.1,4449.7,4252.8,3658.0,0.0000,-396.33,-121.11,-87.953,-47.926,-82.496,-587.69,0.0000,-1050.6,-1520.5,-745.15,-1186.1
1465.000000000,94.359,2181.7,2251.5,1451.4,320.13,3010.7,968.25,5.0184,5656.9,2733.8,3367.3,2069.0,0.0000,-6533.2,-6832.8,-1156.7,-1994.8,-1739.7,-15325.,-99.911,-19012.,-6083.3,-3960.4,-2261.1,71.659,2552.8,2327.7,1500.2,354.61,3162.6,1686.6,0.0000,6719.4,4449.7,4252.8,3658.0,0.0000,-395.01,-120.69,-87.603,-47.772,-82.056,-587.69,0.0000,-1050.6,-1520.4,-745.14,-1186.0
1466.000000000,93.994,2174.7,2244.7,1445.2,319.15,2997.3,968.25,5.0137,5648.6,2733.7,3367.2,2069.1,0.0000,-6530.4,-6830.9,-1155.1,-1994.1,-1736.8,-15324.,-99.877,-19010.,-6082.9,-3960.0,-2260.6,71.446,2545.2,2320.8,1494.0,353.53,3148.8,1686.6,0.0000,6711.1,4449.7,4252.8,3658.0,0.0000,-393.80,-120.30,-87.273,-47.630,-81.634,-587.69,0.0000,-1050.5,-1520.4,-745.13,-1185.9
1467.000000000,94.127,2168.1,2238.3,1439.1,318.17,2984.6,968.25,4.0087,5640.6,2733.7,3367.2,2069.1,0.0000,-6527.3,-6829.0,-1153.6,-1993.4,-1733.9,-15322.,-99.843,-19008.,-6082.5,-3959.6,-2260.1,71.240,2537.9,2314.1,1487.9,352.48,3135.3,1686.6,0.0000,6702.9,4449.7,4252.8,3658.0,0.0000,-392.62,-119.93,-86.952,-47.494,-81.217,-587.69,0.0000,-1050.4,-1520.3,-745.11,-1185.8
1468.000000000,93.618,2161.8,2232.0,1433.0,317.26,2971.6,968.25,3.2006,5633.2,2734.0,3367.2,2069.3,0.0000,-6524.1,-6827.1,-1152.0,-1992.6,-1730.9,-15321.,-99.809,-19006.,-6082.1,-3959.1,-2259.6,71.078,2532.1,2308.9,1482.6,351.64,3123.4,1686.6,0.0000,6695.7,4449.7,4252.8,3658.0,0.0000,-391.68,-119.62,-86.681,-47.386,-80.842,-587.69,0.0000,-1050.3,-1520.3,-745.10,-1185.7
1469.000000000,93.416,2156.2,2226.1,1427.2,316.45,2959.0,968.25,4.8038,5625.3,2734.6,3367.1,2069.4,0.0000,-6520.8,-6825.2,-1150.4,-1991.9,-1727.9,-15319.,-99.775,-19004.,-6081.8,-3958.7,-2259.1,70.908,2526.1,2303.3,1477.2,350.77,3111.2,1686.6,0.0000,6688.3,4449.7,4252.8,3658.0,0.0000,-390.69,-119.30,-86.400,-47.272,-80.460,-587.69,0.0000,-1050.3,-1520.2,-745.09,-1185.6
1470.000000000,93.232,2150.5,2220.3,1421.6,315.64,2947.6,968.25,5.1738,5617.8,2734.8,3367.1,2069.5,0.0000,-6517.4,-6823.2,-1148.8,-1991.1,-1724.9,-15317.,-99.741,-19002.,-6081.4,-3958.2,-2258.6,70.719,2519.3,2297.2,1471.4,349.80,3098.4,1686.6,0.0000,6680.5,4449.7,4252.8,3658.0,0.0000,-389.60,-118.95,-86.098,-47.146,-80.062,-587.69,0.0000,-1050.2,-1520.1,-745.08,-1185.5
1471.000000000,93.048,2144.7,2214.5,1416.0,314.77,2937.5,968.25,5.1737,5609.9,2734.6,3367.1,2069.5,0.0000,-6513.9,-6821.2,-1147.2,-1990.3,-1721.9,-15316.,-99.707,-19001.,-6081.0,-3957.8,-2258.1,70.499,2511.5,2290.1,1465.2,348.68,3084.5,1686.6,0.0000,6672.1,4449.7,4252.8,3658.0,0.0000,-388.33,-118.54,-85.763,-46.999,-79.635,-587.69,0.0000,-1050.1,-1520.1,-745.07,-1185.4
1472.000000000,92.846,2138.6,2208.0,1410.5,313.79,2924.9,968.24,5.1786,5602.2,2734.8,3367.0,2069.6,0.0000,-6510.2,-6819.2,-1145.5,-1989.6,-1718.8,-15314.,-99.673,-18999.,-6080.6,-3957.4,-2257.6,70.260,2503.0,2282.3,1458.5,347.47,3070.0,1686.6,0.0000,6663.4,4449.7,4252.8,3658.0,0.0000,-386.96,-118.10,-85.406,-46.840,-79.191,-587.69,0.0000,-1050.1,-1520.0,-745.05,-1185.3
1473.000000000,92.626,2132.0,2201.0,1404.7,312.78,2912.0,968.21,3.9717,5594.9,2734.8,3367.0,2069.6,0.0000,-6506.3,-6817.1,-1143.9,-1988.8,-1715.8,-15312.,-99.639,-18997.,-6080.2,-3956.9,-2257.1,70.021,2494.5,2274.5,1451.9,346.26,3055.5,1686.6,0.0000,6654.6,4449.7,4252.8,3658.0,0.0000,-385.58,-117.66,-85.050,-46.681,-78.748,-587.69,0.0000,-1050.0,-1519.9,-745.04,-1185.3
1474.000000000,92.395,2125.1,2193.9,1398.8,311.75,2899.2,968.21,3.3678,5587.8,2734.8,3367.0,2069.7,0.0000,-6502.3,-6814.9,-1142.2,-1988.0,-1712.6,-15311.,-99.605,-18995.,-6079.8,-3956.5,-2256.6,69.782,2485.9,2266.8,1445.3,345.05,3041.0,1686.6,0.0000,6645.8,4449.7,4252.8,3658.0,0.0000,-384.21,-117.22,-84.693,-46.521,-78.304,-587.69,0.0000,-1049.9,-1519.9,-745.03,-1185.2
1475.000000000,92.156,2118.6,2187.1,1392.8,310.81,2886.5,968.21,3.3684,5580.5,2734.9,3366.9,2069.8,0.0000,-6498.2,-6812.8,-1140.6,-1987.1,-1709.5,-15309.,-99.572,-18993.,-6079.4,-3956.0,-2256.1,69.614,2479.9,2261.3,1440.8,344.20,3031.3,1686.6,0.0000,6639.9,4449.7,4252.8,3658.0,0.0000,-383.22,-116.90,-84.447,-46.409,-77.987,-587.69,0.0000,-1049.8,-1519.8,-745.02,-1185.1
1476.000000000,91.955,2113.2,2181.4,1387.1,309.97,2874.3,968.20,3.0113,5573.1,2735.2,3366.9,2069.9,0.0000,-6494.0,-6810.6,-1138.9,-1986.3,-1706.3,-15308.,-99.538,-18991.,-6079.1,-3955.6,-2255.6,69.533,2477.1,2258.7,1437.1,343.77,3022.7,1686.6,0.0000,6634.7,4449.7,4252.8,3658.0,0.0000,-382.71,-116.72,-84.272,-46.355,-77.699,-587.69,0.0000,-1049.8,-1519.8,-745.00,-1185.0
1477.000000000,91.873,2111.2,2178.6,1382.0,309.74,2863.2,968.17,2.8250,5565.9,2735.5,3366.9,2070.0,0.0000,-6490.0,-6808.6,-1137.3,-1985.5,-1703.2,-15306.,-99.505,-18989.,-6078.7,-3955.1,-2255.1,206.18,2524.2,2328.8,1448.2,350.09,3028.4,1686.6,13.234,6639.3,4452.1,4256.3,3660.7,0.0000,-384.52,-118.51,-84.442,-46.605,-77.597,-587.69,-0.60423,-1049.8,-1519.7,-745.01,-1184.9
1478.000000000,92.084,2113.7,2178.6,1377.9,309.96,2853.0,968.17,2.8255,5559.1,2735.5,3366.9,2070.1,0.0000,-6486.4,-6806.8,-1135.6,-1984.8,-1700.1,-15304.,-99.473,-18987.,-6078.3,-3954.7,-2254.6,69.746,2484.7,2265.6,1431.9,344.66,3006.5,1686.6,0.0000,6624.9,4449.7,4252.8,3658.0,0.0000,-383.76,-117.01,-84.184,-46.497,-77.148,-587.69,0.0000,-1049.7,-1519.6,-744.98,-1184.8
1479.000000000,92.031,2115.0,2179.2,1374.5,310.08,2843.3,968.16,2.8261,5552.2,2735.4,3366.9,2070.1,0.0000,-6483.1,-6805.2,-1134.0,-1984.1,-1697.0,-15303.,-99.440,-18985.,-6077.9,-3954.3,-2254.0,201.14,2595.1,2353.6,1465.6,360.67,3025.6,1686.6,80.686,6644.6,4459.9,4263.0,3666.8,0.0000,-385.94,-119.23,-84.454,-46.836,-77.221,-587.69,-3.6840,-1049.9,-1519.6,-745.02,-1184.8
1480.000000000,92.275,2118.7,2181.7,1371.2,310.94,2834.2,968.01,3.0949,5545.6,2735.5,3366.9,2070.2,0.0000,-6480.3,-6803.8,-1132.5,-1983.4,-1693.9,-15301.,-99.408,-18983.,-6077.5,-3953.8,-2253.5,70.129,2498.3,2278.0,1430.0,346.38,2997.4,1686.6,0.0000,6619.2,4449.7,4252.8,3658.0,0.0000,-385.77,-117.59,-84.300,-46.753,-76.783,-587.69,0.0000,-1049.5,-1519.5,-744.95,-1184.6
1481.000000000,92.339,2119.6,2183.0,1368.7,310.93,2825.0,968.00,4.8006,5539.0,2735.5,3366.9,2070.3,0.0000,-6477.6,-6802.6,-1130.9,-1982.7,-1690.8,-15299.,-99.375,-18981.,-6077.1,-3953.4,-2253.0,70.032,2494.9,2274.9,1424.6,345.85,2984.5,1686.6,0.0000,6611.4,4449.7,4252.8,3658.0,0.0000,-385.19,-117.40,-84.060,-46.688,-76.383,-587.69,0.0000,-1049.5,-1519.5,-744.94,-1184.5
1482.000000000,92.352,2118.0,2181.3,1365.5,310.92,2815.1,968.00,4.5463,5532.5,2735.6,3366.9,2070.3,0.0000,-6474.8,-6801.3,-1129.4,-1982.0,-1687.7,-15298.,-99.342,-18979.,-6076.7,-3952.9,-2252.5,69.887,2489.7,2270.2,1418.9,345.08,2971.1,1686.6,0.0000,6603.3,4449.7,4252.8,3658.0,0.0000,-384.34,-117.13,-83.782,-46.591,-75.972,-587.69,0.0000,-1049.4,-1519.4,-744.93,-1184.4
1483.000000000,92.305,2114.8,2178.5,1362.0,310.42,2804.6,967.99,2.9865,5526.4,2735.6,3367.0,2070.4,0.0000,-6471.9,-6799.9,-1127.8,-1981.3,-1684.6,-15296.,-99.309,-18977.,-6076.4,-3952.5,-2252.0,69.712,2483.4,2264.5,1412.8,344.18,2957.5,1686.6,0.0000,6595.1,4449.7,4252.8,3658.0,0.0000,-383.32,-116.81,-83.480,-46.475,-75.553,-587.69,0.0000,-1049.3,-1519.3,-744.92,-1184.3
1484.000000000,92.280,2110.8,2174.8,1357.4,309.74,2794.0,967.99,2.9874,5520.4,2735.6,3367.0,2070.5,0.0000,-6468.9,-6798.4,-1126.2,-1980.6,-1681.4,-15294.,-99.275,-18975.,-6076.0,-3952.0,-2251.5,69.543,2477.4,2259.0,1407.1,343.31,2944.6,1686.6,0.0000,6587.3,4449.7,4252.8,3658.0,0.0000,-382.34,-116.50,-83.192,-46.362,-75.154,-587.69,0.0000,-1049.3,-1519.3,-744.90,-1184.2
1485.000000000,92.164,2106.5,2170.5,1352.6,308.94,2783.8,967.83,2.9904,5514.9,2735.7,3367.0,2070.6,0.0000,-6465.8,-6796.9,-1124.6,-1979.8,-1678.2,-15292.,-99.242,-18973.,-6075.6,-3951.6,-2251.0,69.357,2470.8,2253.0,1401.3,342.35,2931.4,1686.6,0.0000,6579.3,4449.7,4252.8,3658.0,0.0000,-381.27,-116.16,-82.889,-46.238,-74.748,-587.69,0.0000,-1049.2,-1519.2,-744.89,-1184.1
1486.000000000,91.985,2101.7,2165.6,1347.6,308.09,2773.4,967.83,3.9480,5509.0,2735.6,3366.9,2070.6,0.0000,-6462.4,-6795.3,-1123.0,-1979.1,-1675.0,-15291.,-99.208,-18971.,-6075.2,-3951.2,-2250.5,69.141,2463.1,2246.0,1395.0,341.25,2917.6,1686.6,0.0000,6570.9,4449.7,4252.8,3658.0,0.0000,-380.03,-115.76,-82.558,-46.094,-74.323,-587.69,0.0000,-1049.1,-1519.2,-744.88,-1184.0
1487.000000000,91.786,2096.7,2160.4,1342.3,307.28,2763.0,967.83,3.6432,5503.5,2735.6,3366.9,2070.8,0.0000,-6459.0,-6793.6,-1121.3,-1978.3,-1671.7,-15289.,-99.175,-18969.,-6074.8,-3950.7,-2250.0,68.963,2456.8,2240.2,1389.4,340.34,2905.1,1686.6,0.0000,6563.4,4449.7,4252.8,3658.0,0.0000,-378.99,-115.43,-82.270,-45.975,-73.936,-587.69,0.0000,-1049.0,-1519.1,-744.87,-1183.9
1488.000000000,91.600,2091.6,2155.1,1337.1,306.42,2752.3,967.83,2.6058,5497.4,2735.6,3366.9,2070.9,0.0000,-6455.3,-6791.9,-1119.7,-1977.5,-1668.4,-15287.,-99.141,-18967.,-6074.4,-3950.3,-2249.5,68.783,2450.3,2234.3,1383.9,339.42,2892.8,1686.6,0.0000,6555.9,4449.7,4252.8,3658.0,0.0000,-377.94,-115.10,-81.981,-45.855,-73.551,-587.69,0.0000,-1049.0,-1519.0,-744.85,-1183.8
1489.000000000,91.412,2086.7,2150.0,1331.9,305.63,2741.3,967.83,2.6064,5490.8,2735.6,3366.9,2071.0,0.0000,-6451.6,-6790.1,-1118.0,-1976.7,-1665.1,-15286.,-99.108,-18965.,-6074.0,-3949.8,-2249.0,68.642,2445.4,2229.8,1379.1,338.69,2881.8,1686.6,0.0000,6549.2,4449.7,4252.8,3658.0,0.0000,-377.11,-114.83,-81.736,-45.762,-73.201,-587.69,0.0000,-1048.9,-1519.0,-744.84,-1183.7
1490.000000000,91.209,2082.4,2145.2,1326.8,304.90,2730.0,967.83,2.6069,5483.9,2735.7,3366.9,2071.1,0.0000,-6447.8,-6788.4,-1116.3,-1975.9,-1661.7,-15284.,-99.074,-18963.,-6073.6,-3949.4,-2248.5,68.467,2439.1,2224.0,1373.7,337.79,2869.8,1686.6,0.0000,6542.0,4449.7,4252.8,3658.0,0.0000,-376.09,-114.50,-81.456,-45.644,-72.828,-587.69,0.0000,-1048.8,-1518.9,-744.83,-1183.6
1491.000000000,91.031,2077.5,2140.5,1321.7,304.12,2718.6,967.83,2.6075,5477.2,2735.6,3366.8,2071.2,0.0000,-6443.9,-6786.6,-1114.6,-1975.1,-1658.4,-15282.,-99.041,-18961.,-6073.3,-3948.9,-2248.0,68.275,2432.3,2217.8,1368.1,336.81,2857.5,1686.6,0.0000,6534.5,4449.7,4252.8,3658.0,0.0000,-374.97,-114.14,-81.160,-45.517,-72.443,-587.69,0.0000,-1048.8,-1518.9,-744.82,-1183.5
1492.000000000,90.851,2072.2,2135.0,1316.6,303.31,2707.2,967.83,2.6080,5470.3,2735.6,3366.7,2071.3,0.0000,-6439.9,-6784.7,-1112.8,-1974.3,-1655.1,-15280.,-99.008,-18959.,-6072.9,-3948.5,-2247.5,68.072,2425.0,2211.2,1362.4,335.78,2844.8,1686.6,0.0000,6526.9,4449.7,4252.8,3658.0,0.0000,-373.79,-113.77,-80.853,-45.381,-72.051,-587.69,0.0000,-1048.7,-1518.8,-744.80,-1183.4
1493.000000000,90.661,2066.7,2129.4,1311.5,302.44,2695.9,967.83,2.6086,5463.2,2735.6,3366.7,2071.4,0.0000,-6435.7,-6782.9,-1111.1,-1973.5,-1651.7,-15279.,-98.974,-18957.,-6072.5,-3948.1,-2247.0,67.857,2417.4,2204.2,1356.4,334.70,2831.8,1686.6,0.0000,6519.0,4449.7,4252.8,3658.0,0.0000,-372.55,-113.37,-80.533,-45.238,-71.650,-587.69,0.0000,-1048.6,-1518.7,-744.79,-1183.3
1494.000000000,90.455,2060.8,2123.4,1306.6,301.52,2684.4,967.83,3.1341,5456.2,2735.7,3366.7,2071.5,0.0000,-6431.5,-6780.9,-1109.4,-1972.6,-1648.3,-15277.,-98.941,-18955.,-6072.1,-3947.6,-2246.5,67.637,2409.5,2197.1,1350.4,333.58,2818.7,1686.6,0.0000,6511.1,4449.7,4252.8,3658.0,0.0000,-371.27,-112.96,-80.208,-45.092,-71.245,-587.69,0.0000,-1048.5,-1518.7,-744.78,-1183.2
1495.000000000,90.246,2054.7,2117.4,1301.3,300.60,2672.8,967.83,4.0384,5449.3,2735.7,3366.6,2071.6,0.0000,-6427.1,-6778.9,-1107.6,-1971.8,-1644.9,-15275.,-98.908,-18953.,-6071.7,-3947.2,-2246.0,67.445,2402.7,2190.9,1344.9,332.61,2806.5,1686.6,0.0000,6503.7,4449.7,4252.8,3658.0,0.0000,-370.15,-112.60,-79.914,-44.963,-70.865,-587.69,0.0000,-1048.5,-1518.6,-744.77,-1183.1
1496.000000000,90.059,2049.0,2111.5,1296.0,299.61,2661.2,967.84,4.0388,5442.3,2735.8,3366.6,2071.7,0.0000,-6422.6,-6776.9,-1105.8,-1970.9,-1641.5,-15274.,-98.875,-18951.,-6071.3,-3946.7,-2245.5,67.258,2396.0,2184.8,1339.4,331.66,2794.5,1686.6,0.0000,6496.4,4449.7,4252.8,3658.0,0.0000,-369.05,-112.25,-79.626,-44.839,-70.491,-587.69,0.0000,-1048.4,-1518.6,-744.75,-1183.0
1497.000000000,89.859,2043.4,2105.6,1290.8,298.79,2649.8,967.84,4.0392,5435.4,2735.8,3366.6,2071.8,0.0000,-6418.1,-6774.8,-1104.1,-1970.1,-1638.1,-15272.,-98.842,-18949.,-6070.9,-3946.3,-2245.0,67.066,2389.2,2178.5,1334.0,330.68,2782.6,1686.6,0.0000,6489.3,4449.7,4252.8,3658.0,0.0000,-367.93,-111.89,-79.337,-44.711,-70.120,-587.69,0.0000,-1048.3,-1518.5,-744.74,-1183.0
1498.000000000,89.661,2037.5,2099.6,1285.8,297.92,2638.6,967.84,2.2699,5428.6,2735.9,3366.5,2071.9,0.0000,-6413.5,-6772.7,-1102.3,-1969.2,-1634.6,-15270.,-98.808,-18946.,-6070.5,-3945.8,-2244.5,66.843,2381.2,2171.3,1328.1,329.55,2769.6,1686.6,0.0000,6481.4,4449.7,4252.8,3658.0,0.0000,-366.63,-111.48,-79.011,-44.562,-69.719,-587.69,0.0000,-1048.2,-1518.4,-744.73,-1182.9
1499.000000000,89.577,2031.3,2093.0,1280.6,297.00,2627.6,967.83,2.2248,5422.0,2735.8,3366.5,2072.0,0.0000,-6408.7,-6770.5,-1100.5,-1968.3,-1631.2,-15268.,-98.775,-18944.,-6070.1,-3945.4,-2244.0,66.611,2373.0,2163.8,1322.0,328.39,2756.3,1686.6,0.0000,6473.4,4449.7,4252.8,3658.0,0.0000,-365.29,-111.05,-78.678,-44.408,-69.312,-587.69,0.0000,-1048.2,-1518.4,-744.71,-1182.8
1500.000000000,89.387,2024.9,2086.8,1275.3,296.08,2616.3,967.83,2.2253,5415.0,2735.8,3366.5,2072.0,0.0000,-6403.9,-6768.2,-1098.7,-1967.4,-1627.7,-15267.,-98.742,-18942.,-6069.7,-3944.9,-2243.5,66.382,2364.8,2156.3,1315.9,327.23,2743.1,1686.6,0.0000,6465.4,4449.7,4252.8,3658.0,0.0000,-363.96,-110.62,-78.346,-44.255,-68.907,-587.69,0.0000,-1048.1,-1518.3,-744.70,-1182.7
1501.000000000,89.162,2018.5,2080.3,1269.9,295.06,2604.7,967.83,2.2258,5408.1,2735.9,3366.4,2072.1,0.0000,-6399.0,-6765.9,-1096.8,-1966.5,-1624.2,-15265.,-98.709,-18940.,-6069.3,-3944.5,-2243.0,66.157,2356.8,2149.0,1309.9,326.10,2730.0,1686.6,0.0000,6457.5,4449.7,4252.8,3658.0,0.0000,-362.64,-110.20,-78.019,-44.105,-68.505,-587.69,0.0000,-1048.0,-1518.3,-744.69,-1182.6
1502.000000000,88.867,2011.9,2074.0,1264.4,294.07,2592.9,967.83,2.2263,5401.1,2736.0,3366.5,2072.1,0.0000,-6394.0,-6763.6,-1095.0,-1965.6,-1620.7,-15263.,-98.676,-18938.,-6068.9,-3944.0,-2242.5,65.945,2349.3,2142.1,1304.1,325.02,2717.4,1686.6,0.0000,6449.8,4449.7,4252.8,3658.0,0.0000,-361.40,-109.80,-77.706,-43.963,-68.115,-587.69,0.0000,-1048.0,-1518.2,-744.68,-1182.5
1503.000000000,88.497,2005.6,2067.4,1258.9,293.10,2581.5,967.83,2.2269,5394.1,2736.1,3366.4,2072.2,0.0000,-6388.9,-6761.2,-1093.1,-1964.7,-1617.1,-15261.,-98.643,-18936.,-6068.5,-3943.6,-2242.0,65.717,2341.1,2134.7,1298.0,323.87,2704.3,1686.6,0.0000,6441.9,4449.7,4252.8,3658.0,0.0000,-360.07,-109.38,-77.377,-43.811,-67.714,-587.69,0.0000,-1047.9,-1518.1,-744.66,-1182.4
1504.000000000,88.227,1999.1,2060.8,1253.4,292.14,2569.9,967.83,2.2274,5387.2,2736.1,3366.4,2072.2,0.0000,-6383.8,-6758.8,-1091.3,-1963.7,-1613.5,-15260.,-98.610,-18934.,-6068.2,-3943.2,-2241.5,65.475,2332.5,2126.8,1291.8,322.65,2690.8,1686.6,0.0000,6433.7,4449.7,4252.8,3658.0,0.0000,-358.66,-108.93,-77.033,-43.650,-67.301,-587.69,0.0000,-1047.8,-1518.1,-744.65,-1182.3
1505.000000000,87.973,1992.3,2054.2,1248.0,291.13,2558.2,967.83,2.2280,5380.4,2736.1,3366.4,2072.3,0.0000,-6378.7,-6756.4,-1089.4,-1962.8,-1610.0,-15258.,-98.577,-18932.,-6067.8,-3942.7,-2241.0,65.251,2324.5,2119.6,1285.8,321.53,2677.9,1686.6,0.0000,6425.9,4449.7,4252.8,3658.0,0.0000,-357.35,-108.51,-76.709,-43.501,-66.904,-587.69,0.0000,-1047.7,-1518.0,-744.64,-1182.2
1506.000000000,87.583,1997.1,2057.6,1242.8,292.10,2548.0,967.83,2.2285,5373.6,2736.2,3366.4,2072.4,0.0000,-6374.2,-6754.4,-1087.6,-1961.9,-1606.4,-15256.,-98.546,-18930.,-6067.4,-3942.3,-2240.5,134.49,2445.8,2231.9,1317.4,335.52,2724.7,1686.6,31.729,6455.5,4452.2,4255.4,3660.4,0.0000,-369.48,-113.02,-78.723,-44.999,-67.957,-587.69,-1.4487,-1047.8,-1517.9,-744.64,-1182.1
1507.000000000,88.473,2024.2,2079.8,1240.2,296.38,2542.2,967.83,2.2290,5368.1,2736.3,3366.4,2072.4,0.0000,-6371.9,-6753.7,-1086.0,-1961.3,-1603.0,-15254.,-98.516,-18927.,-6067.0,-3941.8,-2240.0,68.280,2432.4,2218.0,1314.4,336.61,2716.8,1686.6,0.0000,6449.1,4449.9,4253.1,3658.2,0.0000,-373.82,-113.49,-79.192,-45.524,-67.751,-587.69,0.0000,-1047.7,-1517.9,-744.61,-1182.0
1508.000000000,89.217,2045.4,2101.1,1242.3,298.59,2538.9,967.82,2.2296,5362.9,2736.2,3366.4,2072.5,0.0000,-6370.8,-6754.0,-1084.5,-1960.9,-1599.6,-15253.,-98.485,-18925.,-6066.6,-3941.4,-2239.5,68.411,2437.1,2222.2,1310.9,337.08,2706.5,1686.6,0.0000,6442.8,4449.9,4253.0,3658.2,0.0000,-374.49,-113.70,-79.138,-45.611,-67.423,-587.69,0.0000,-1047.6,-1517.8,-744.60,-1181.9
1509.000000000,89.913,2054.9,2110.6,1244.1,301.18,2535.0,967.79,2.2301,5358.4,2736.2,3366.4,2072.6,0.0000,-6370.1,-6754.2,-1083.0,-1960.4,-1596.5,-15251.,-98.453,-18923.,-6066.2,-3941.0,-2239.0,68.403,2436.8,2222.0,1306.8,336.71,2696.1,1686.6,0.0000,6436.5,4449.8,4252.9,3658.1,0.0000,-374.41,-113.68,-78.992,-45.604,-67.097,-587.69,0.0000,-1047.6,-1517.8,-744.59,-1181.8
1510.000000000,90.458,2057.6,2114.4,1243.9,302.16,2528.6,967.79,2.2306,5353.3,2736.3,3366.4,2072.7,0.0000,-6369.3,-6754.2,-1081.5,-1959.9,-1593.2,-15249.,-98.421,-18921.,-6065.8,-3940.5,-2238.5,68.283,2432.6,2218.1,1301.5,335.94,2684.1,1686.6,0.0000,6429.2,4449.7,4252.9,3658.1,0.0000,-373.71,-113.46,-78.751,-45.524,-66.730,-587.69,0.0000,-1047.5,-1517.7,-744.57,-1181.7
1511.000000000,90.548,2057.2,2114.3,1242.2,301.95,2520.8,967.79,2.2311,5347.6,2736.4,3366.4,2072.8,0.0000,-6368.2,-6754.0,-1079.9,-1959.3,-1589.9,-15247.,-98.389,-18919.,-6065.4,-3940.1,-2238.0,68.111,2426.4,2212.5,1295.9,334.94,2671.7,1686.6,0.0000,6421.6,4449.7,4252.8,3658.0,0.0000,-372.73,-113.16,-78.469,-45.408,-66.351,-587.69,0.0000,-1047.4,-1517.6,-744.56,-1181.6
1512.000000000,90.626,2055.4,2112.7,1239.9,301.50,2512.7,967.79,2.2316,5342.8,2736.4,3366.3,2072.9,0.0000,-6366.8,-6753.7,-1078.5,-1958.7,-1586.6,-15245.,-98.356,-18917.,-6065.1,-3939.6,-2237.5,68.068,2424.9,2211.1,1292.9,334.62,2664.4,1686.6,0.0000,6417.2,4449.8,4252.8,3658.0,0.0000,-372.47,-113.08,-78.339,-45.379,-66.104,-587.69,0.0000,-1047.3,-1517.6,-744.55,-1181.5
1513.000000000,90.468,2053.2,2112.0,1237.1,301.02,2503.2,967.79,2.2322,5337.9,2736.5,3366.3,2073.0,0.0000,-6365.3,-6753.1,-1076.9,-1958.1,-1583.2,-15244.,-98.324,-18915.,-6064.7,-3939.2,-2237.1,67.870,2417.8,2204.7,1287.5,333.62,2652.5,1686.6,0.0000,6410.0,4449.7,4252.8,3658.0,0.0000,-371.34,-112.74,-78.046,-45.247,-65.738,-587.69,0.0000,-1047.3,-1517.5,-744.53,-1181.4
1514.000000000,90.102,2050.9,2110.6,1233.0,300.20,2494.9,967.79,2.2327,5335.2,2736.5,3366.3,2073.0,0.0000,-6363.6,-6752.4,-1075.3,-1957.4,-1579.7,-15242.,-98.291,-18913.,-6064.3,-3938.8,-2236.6,67.648,2409.9,2197.4,1281.7,332.47,2640.1,1686.6,0.0000,6402.5,4449.7,4252.8,3658.0,0.0000,-370.09,-112.35,-77.732,-45.099,-65.362,-587.69,0.0000,-1047.2,-1517.5,-744.52,-1181.3
1515.000000000,89.835,2046.4,2106.0,1229.4,299.36,2488.7,967.79,2.2332,5333.5,2736.5,3366.3,2073.1,0.0000,-6361.7,-6751.6,-1073.7,-1956.7,-1576.3,-15240.,-98.259,-18911.,-6063.9,-3938.3,-2236.1,67.405,2401.3,2189.6,1275.8,331.25,2627.4,1686.6,0.0000,6394.8,4449.7,4252.8,3658.0,0.0000,-368.72,-111.93,-77.399,-44.937,-64.976,-587.69,0.0000,-1047.1,-1517.4,-744.51,-1181.2
1516.000000000,89.629,2040.5,2100.2,1225.5,298.37,2482.4,967.80,2.2337,5330.5,2736.6,3366.4,2073.2,0.0000,-6359.3,-6750.5,-1072.0,-1956.0,-1572.8,-15238.,-98.226,-18909.,-6063.5,-3937.9,-2235.6,67.149,2392.1,2181.2,1269.7,329.96,2614.4,1686.6,0.0000,6386.9,4449.7,4252.8,3658.0,0.0000,-367.27,-111.48,-77.054,-44.766,-64.584,-587.69,0.0000,-1047.1,-1517.3,-744.50,-1181.1
1517.000000000,89.387,2035.9,2093.8,1220.9,297.33,2474.6,967.80,2.2342,5326.0,2736.6,3366.4,2073.3,0.0000,-6356.6,-6749.3,-1070.4,-1955.3,-1569.3,-15236.,-98.194,-18906.,-6063.1,-3937.5,-2235.1,66.928,2384.3,2174.0,1264.1,328.85,2602.6,1686.6,0.0000,6379.8,4449.7,4252.8,3658.0,0.0000,-366.01,-111.08,-76.748,-44.618,-64.223,-587.69,0.0000,-1047.0,-1517.3,-744.48,-1181.0
1518.000000000,89.122,2030.4,2088.4,1216.3,296.33,2464.9,967.80,2.2347,5320.7,2736.6,3366.4,2073.4,0.0000,-6353.7,-6748.0,-1068.7,-1954.5,-1565.7,-15235.,-98.161,-18904.,-6062.8,-3937.1,-2234.6,66.716,2376.7,2167.2,1258.9,327.79,2591.2,1686.6,0.0000,6373.0,4449.7,4252.8,3658.0,0.0000,-364.81,-110.71,-76.453,-44.478,-63.873,-587.69,0.0000,-1046.9,-1517.2,-744.47,-1181.0
1519.000000000,88.655,2024.4,2082.7,1211.7,295.25,2454.4,967.80,2.2352,5314.9,2736.7,3366.4,2073.5,0.0000,-6350.5,-6746.6,-1066.9,-1953.7,-1562.2,-15233.,-98.128,-18902.,-6062.4,-3936.6,-2234.1,66.477,2368.2,2159.4,1253.2,326.60,2579.1,1686.6,0.0000,6365.7,4449.7,4252.8,3658.0,0.0000,-363.44,-110.28,-76.131,-44.318,-63.504,-587.69,0.0000,-1046.9,-1517.1,-744.46,-1180.9
1520.000000000,88.419,2018.3,2076.9,1206.6,294.19,2443.6,967.80,2.2444,5308.7,2736.7,3366.4,2073.6,0.0000,-6347.1,-6745.2,-1065.2,-1953.0,-1558.6,-15231.,-98.096,-18900.,-6062.0,-3936.2,-2233.6,66.212,2358.8,2150.8,1247.1,325.27,2566.3,1686.6,0.0000,6357.9,4449.7,4252.8,3658.0,0.0000,-361.93,-109.81,-75.782,-44.141,-63.117,-587.69,0.0000,-1046.8,-1517.1,-744.44,-1180.8
1521.000000000,88.172,2011.3,2071.0,1201.4,293.09,2433.0,967.80,2.2641,5302.4,2736.8,3366.4,2073.7,0.0000,-6343.7,-6743.6,-1063.4,-1952.2,-1555.0,-15229.,-98.063,-18898.,-6061.6,-3935.8,-2233.1,65.946,2349.3,2142.2,1241.0,323.95,2553.4,1686.6,0.0000,6350.1,4449.7,4252.8,3658.0,0.0000,-360.42,-109.34,-75.432,-43.964,-62.729,-587.69,0.0000,-1046.7,-1517.0,-744.43,-1180.7
1522.000000000,87.918,2005.1,2064.1,1196.1,292.01,2422.6,967.80,2.2646,5296.0,2736.8,3366.3,2073.8,0.0000,-6340.1,-6741.9,-1061.6,-1951.3,-1551.4,-15228.,-98.030,-18896.,-6061.2,-3935.4,-2232.6,65.726,2341.5,2135.0,1235.6,322.85,2542.0,1686.6,0.0000,6343.2,4449.7,4252.8,3658.0,0.0000,-359.16,-108.94,-75.132,-43.818,-62.378,-587.69,0.0000,-1046.6,-1517.0,-744.42,-1180.6
1523.000000000,87.679,1999.0,2057.4,1190.7,290.99,2412.5,967.80,2.2651,5290.0,2736.8,3366.3,2073.8,0.0000,-6336.3,-6740.2,-1059.8,-1950.5,-1547.8,-15226.,-97.998,-18894.,-6060.9,-3935.0,-2232.1,65.511,2333.8,2128.0,1230.4,321.77,2530.8,1686.6,0.0000,6336.5,4449.7,4252.8,3658.0,0.0000,-357.92,-108.54,-74.837,-43.674,-62.033,-587.69,0.0000,-1046.6,-1516.9,-744.40,-1180.5
1524.000000000,87.445,1992.7,2050.7,1185.5,290.01,2402.7,967.80,2.2656,5283.6,2736.9,3366.4,2073.9,0.0000,-6332.4,-6738.4,-1058.0,-1949.7,-1544.2,-15224.,-97.965,-18892.,-6060.5,-3934.6,-2231.6,65.298,2326.2,2121.1,1225.2,320.70,2519.7,1686.6,0.0000,6329.7,4449.7,4252.8,3658.0,0.0000,-356.68,-108.15,-74.544,-43.532,-61.690,-587.69,0.0000,-1046.5,-1516.8,-744.39,-1180.4
1525.000000000,87.220,1986.9,2044.3,1180.9,289.16,2392.1,967.80,2.2661,5277.0,2736.9,3366.4,2074.0,0.0000,-6328.4,-6736.5,-1056.2,-1948.8,-1540.5,-15222.,-97.933,-18889.,-6060.1,-3934.2,-2231.1,65.163,2321.4,2116.7,1221.2,320.02,2510.8,1686.6,0.0000,6324.4,4449.7,4252.8,3658.0,0.0000,-355.87,-107.89,-74.333,-43.442,-61.405,-587.69,0.0000,-1046.4,-1516.8,-744.38,-1180.3
1526.000000000,87.006,1981.5,2038.3,1176.2,288.40,2381.7,967.80,2.2665,5270.4,2737.0,3366.4,2074.0,0.0000,-6324.3,-6734.6,-1054.4,-1948.0,-1536.9,-15220.,-97.901,-18887.,-6059.7,-3933.8,-2230.6,64.920,2312.7,2108.8,1215.5,318.80,2498.9,1686.6,0.0000,6317.2,4449.7,4252.8,3658.0,0.0000,-354.46,-107.45,-74.010,-43.280,-61.041,-587.69,0.0000,-1046.4,-1516.7,-744.37,-1180.2
1527.000000000,86.630,1975.3,2031.8,1171.7,287.45,2371.2,967.80,2.2670,5264.3,2737.0,3366.4,2074.1,0.0000,-6320.1,-6732.6,-1052.5,-1947.1,-1533.3,-15218.,-97.868,-18885.,-6059.3,-3933.3,-2230.1,64.652,2303.2,2100.1,1209.5,317.47,2486.2,1686.6,0.0000,6309.5,4449.7,4252.8,3658.0,0.0000,-352.92,-106.96,-73.661,-43.101,-60.660,-587.69,0.0000,-1046.3,-1516.7,-744.35,-1180.1
1528.000000000,86.278,1968.3,2024.9,1167.2,286.48,2360.8,967.80,2.2675,5258.0,2737.0,3366.4,2074.2,0.0000,-6315.8,-6730.5,-1050.7,-1946.2,-1529.6,-15217.,-97.836,-18883.,-6059.0,-3932.9,-2229.6,64.403,2294.3,2092.0,1203.7,316.23,2474.1,1686.6,0.0000,6302.2,4449.7,4252.8,3658.0,0.0000,-351.47,-106.51,-73.333,-42.935,-60.294,-587.69,0.0000,-1046.2,-1516.6,-744.34,-1180.0
1529.000000000,86.046,1961.1,2018.2,1162.2,285.43,2350.3,967.80,2.2680,5251.6,2737.1,3366.3,2074.3,0.0000,-6311.3,-6728.4,-1048.8,-1945.3,-1526.0,-15215.,-97.804,-18881.,-6058.6,-3932.5,-2229.1,64.152,2285.4,2083.9,1198.0,314.98,2462.0,1686.6,0.0000,6294.9,4449.7,4252.8,3658.0,0.0000,-350.02,-106.05,-73.003,-42.768,-59.927,-587.69,0.0000,-1046.2,-1516.5,-744.33,-1179.9
1530.000000000,85.792,1954.1,2012.2,1157.0,284.33,2339.5,967.80,2.2685,5245.1,2737.1,3366.3,2074.3,0.0000,-6306.7,-6726.2,-1046.9,-1944.4,-1522.3,-15213.,-97.771,-18879.,-6058.2,-3932.1,-2228.6,63.894,2276.2,2075.5,1192.1,313.69,2449.6,1686.6,0.0000,6287.4,4449.7,4252.8,3658.0,0.0000,-348.52,-105.58,-72.664,-42.596,-59.555,-587.69,0.0000,-1046.1,-1516.5,-744.31,-1179.8
1531.000000000,85.533,1947.0,2005.2,1151.9,283.20,2328.5,967.80,2.2689,5238.7,2737.2,3366.3,2074.4,0.0000,-6302.0,-6723.8,-1045.0,-1943.5,-1518.6,-15211.,-97.739,-18877.,-6057.8,-3931.7,-2228.1,63.647,2267.4,2067.5,1186.8,312.47,2438.7,1686.6,0.0000,6280.8,4449.7,4252.8,3658.0,0.0000,-347.08,-105.12,-72.353,-42.431,-59.221,-587.69,0.0000,-1046.0,-1516.4,-744.28,-1179.7
1532.000000000,85.282,1939.7,1998.1,1146.8,282.11,2318.0,967.81,2.2770,5232.4,2737.2,3366.3,2074.5,0.0000,-6297.2,-6721.4,-1043.1,-1942.6,-1514.9,-15209.,-97.707,-18874.,-6057.4,-3931.3,-2227.7,63.409,2258.9,2059.7,1181.3,311.28,2426.9,1686.6,0.0000,6273.7,4449.7,4252.8,3658.0,0.0000,-345.69,-104.68,-72.036,-42.273,-58.863,-587.69,0.0000,-1046.0,-1516.4,-744.26,-1179.6
1533.000000000,85.218,1932.7,1991.7,1142.1,281.06,2307.5,967.81,2.2786,5226.4,2737.3,3366.4,2074.6,0.0000,-6292.4,-6719.0,-1041.2,-1941.6,-1511.1,-15208.,-97.675,-18872.,-6057.1,-3930.9,-2227.2,63.194,2251.2,2052.8,1176.1,310.20,2415.8,1686.6,0.0000,6267.0,4449.7,4252.8,3658.0,0.0000,-344.42,-104.28,-71.743,-42.129,-58.524,-587.69,0.0000,-1045.9,-1516.3,-744.23,-1179.5
1534.000000000,85.232,1926.0,1985.8,1137.1,280.08,2297.1,967.81,2.2791,5220.7,2737.3,3366.4,2074.6,0.0000,-6287.5,-6716.5,-1039.3,-1940.7,-1507.4,-15206.,-97.643,-18870.,-6056.7,-3930.5,-2226.7,62.977,2243.5,2045.7,1170.8,309.12,2404.7,1686.6,0.0000,6260.3,4449.7,4252.8,3658.0,0.0000,-343.14,-103.87,-71.449,-41.985,-58.184,-587.69,0.0000,-1045.8,-1516.2,-744.20,-1179.4
1535.000000000,85.005,1919.4,1979.0,1132.1,279.10,2286.7,967.81,2.2795,5214.6,2737.3,3366.4,2074.7,0.0000,-6282.5,-6714.0,-1037.4,-1939.7,-1503.6,-15204.,-97.610,-18868.,-6056.3,-3930.1,-2226.2,62.750,2235.4,2038.3,1165.5,307.98,2393.3,1686.6,0.0000,6253.4,4449.7,4252.8,3658.0,0.0000,-341.80,-103.45,-71.144,-41.833,-57.838,-587.69,0.0000,-1045.7,-1516.2,-744.18,-1179.3
1536.000000000,84.774,1912.8,1972.2,1127.2,278.13,2276.8,967.81,2.2767,5208.4,2737.4,3366.4,2074.8,0.0000,-6277.5,-6711.4,-1035.5,-1938.8,-1499.8,-15202.,-97.578,-18866.,-6055.9,-3929.7,-2225.7,62.525,2227.4,2031.0,1160.1,306.86,2382.0,1686.6,0.0000,6246.6,4449.7,4252.8,3658.0,0.0000,-340.48,-103.03,-70.842,-41.683,-57.494,-587.69,0.0000,-1045.7,-1516.1,-744.15,-1179.2
1537.000000000,84.370,1906.0,1965.4,1122.1,277.14,2266.5,967.81,2.2772,5202.2,2737.5,3366.4,2074.9,0.0000,-6272.3,-6708.9,-1033.5,-1937.8,-1496.1,-15200.,-97.546,-18863.,-6055.6,-3929.3,-2225.2,62.267,2218.2,2022.7,1154.3,305.58,2369.7,1686.6,0.0000,6239.2,4449.7,4252.8,3658.0,0.0000,-338.97,-102.55,-70.506,-41.512,-57.126,-587.69,0.0000,-1045.6,-1516.1,-744.12,-1179.1
1538.000000000,84.130,1898.8,1958.2,1117.1,276.08,2256.2,967.81,2.2777,5195.7,2737.5,3366.4,2075.0,0.0000,-6267.1,-6706.2,-1031.6,-1936.8,-1492.3,-15198.,-97.514,-18861.,-6055.2,-3928.9,-2224.7,62.005,2208.9,2014.1,1148.4,304.27,2357.3,1686.6,0.0000,6231.7,4449.7,4252.8,3658.0,0.0000,-337.44,-102.07,-70.165,-41.337,-56.755,-587.69,0.0000,-1045.5,-1516.0,-744.10,-1179.0
1539.000000000,83.879,1891.3,1950.7,1112.0,275.01,2245.4,967.80,2.2781,5189.2,2737.5,3366.5,2075.1,0.0000,-6261.7,-6703.5,-1029.6,-1935.8,-1488.5,-15197.,-97.482,-18859.,-6054.8,-3928.5,-2224.2,61.746,2199.7,2005.7,1142.5,302.98,2345.0,1686.6,0.0000,6224.2,4449.7,4252.8,3658.0,0.0000,-335.92,-101.59,-69.828,-41.164,-56.387,-587.69,0.0000,-1045.5,-1515.9,-744.07,-1178.9
1540.000000000,83.625,1883.8,1943.2,1106.8,273.83,2234.7,967.77,2.2785,5182.8,2737.6,3366.5,2075.2,0.0000,-6256.2,-6700.8,-1027.6,-1934.8,-1484.7,-15195.,-97.450,-18857.,-6054.4,-3928.1,-2223.7,61.486,2190.4,1997.3,1136.6,301.69,2332.6,1686.6,0.0000,6216.8,4449.7,4252.8,3658.0,0.0000,-334.40,-101.11,-69.490,-40.991,-56.019,-587.69,0.0000,-1045.4,-1515.9,-744.04,-1178.9
1541.000000000,83.364,1876.3,1935.3,1101.5,272.67,2223.9,967.74,2.2790,5176.3,2737.6,3366.5,2075.3,0.0000,-6250.6,-6698.0,-1025.6,-1933.8,-1480.8,-15193.,-97.418,-18854.,-6054.0,-3927.7,-2223.2,61.231,2181.3,1989.0,1130.8,300.42,2320.4,1686.6,0.0000,6209.4,4449.7,4252.8,3658.0,0.0000,-332.91,-100.63,-69.156,-40.821,-55.654,-587.69,0.0000,-1045.3,-1515.8,-744.02,-1178.8
1542.000000000,83.105,1868.7,1927.6,1096.2,271.57,2213.3,967.74,2.2794,5169.9,2737.6,3366.6,2075.4,0.0000,-6244.9,-6695.1,-1023.6,-1932.8,-1476.9,-15191.,-97.386,-18852.,-6053.7,-3927.3,-2222.7,60.972,2172.1,1980.6,1124.9,299.13,2308.1,1686.6,0.0000,6202.0,4449.7,4252.8,3658.0,0.0000,-331.39,-100.15,-68.820,-40.648,-55.288,-587.69,0.0000,-1045.3,-1515.8,-743.99,-1178.7
1543.000000000,82.846,1861.4,1919.8,1090.8,270.46,2202.6,967.74,2.2798,5163.6,2737.7,3366.6,2075.4,0.0000,-6239.0,-6692.2,-1021.6,-1931.8,-1473.1,-15189.,-97.354,-18850.,-6053.3,-3926.9,-2222.2,60.717,2163.0,1972.3,1119.1,297.86,2295.9,1686.6,0.0000,6194.6,4449.7,4252.8,3658.0,0.0000,-329.89,-99.677,-68.486,-40.478,-54.924,-587.69,0.0000,-1045.2,-1515.7,-743.96,-1178.6
1544.000000000,82.587,1854.0,1912.1,1085.5,269.38,2191.8,967.74,2.2803,5157.1,2737.7,3366.6,2075.5,0.0000,-6233.1,-6689.3,-1019.6,-1930.7,-1469.2,-15187.,-97.322,-18848.,-6052.9,-3926.5,-2221.8,60.491,2155.0,1965.0,1113.7,296.73,2284.4,1686.6,0.0000,6187.6,4449.7,4252.8,3658.0,0.0000,-328.54,-99.250,-68.181,-40.327,-54.577,-587.69,0.0000,-1045.1,-1515.6,-743.94,-1178.5
1545.000000000,82.344,1847.0,1904.9,1080.2,268.33,2181.2,967.75,2.2807,5150.6,2737.8,3366.6,2075.6,0.0000,-6227.1,-6686.3,-1017.6,-1929.7,-1465.2,-15185.,-97.290,-18846.,-6052.5,-3926.1,-2221.3,60.264,2146.9,1957.6,1108.3,295.59,2273.0,1686.6,0.0000,6180.7,4449.7,4252.8,3658.0,0.0000,-327.19,-98.821,-67.877,-40.176,-54.234,-587.69,0.0000,-1045.1,-1515.6,-743.91,-1178.4
1546.000000000,82.106,1840.5,1897.7,1075.0,267.31,2170.5,967.75,2.2811,5144.4,2737.8,3366.6,2075.7,0.0000,-6221.1,-6683.4,-1015.5,-1928.7,-1461.3,-15184.,-97.258,-18843.,-6052.2,-3925.7,-2220.8,60.035,2138.7,1950.1,1103.0,294.45,2261.6,1686.6,0.0000,6173.8,4449.7,4252.8,3658.0,0.0000,-325.83,-98.388,-67.571,-40.023,-53.891,-587.69,0.0000,-1045.0,-1515.5,-743.88,-1178.3
1547.000000000,81.903,1833.7,1891.2,1069.8,266.31,2159.8,967.75,2.2767,5137.8,2737.9,3366.7,2075.8,0.0000,-6215.0,-6680.5,-1013.5,-1927.6,-1457.4,-15182.,-97.226,-18841.,-6051.8,-3925.3,-2220.3,59.789,2130.0,1942.2,1097.3,293.23,2249.7,1686.6,0.0000,6166.7,4449.7,4252.8,3658.0,0.0000,-324.39,-97.929,-67.249,-39.860,-53.537,-587.69,0.0000,-1044.9,-1515.4,-743.85,-1178.2
1548.000000000,81.754,1826.6,1884.0,1064.6,265.30,2149.0,967.75,2.2760,5131.2,2737.9,3366.7,2075.9,0.0000,-6208.9,-6677.6,-1011.5,-1926.6,-1453.4,-15180.,-97.194,-18839.,-6051.4,-3924.9,-2219.8,59.545,2121.2,1934.2,1091.7,292.01,2237.8,1686.6,0.0000,6159.5,4449.7,4252.8,3658.0,0.0000,-322.94,-97.471,-66.928,-39.696,-53.184,-587.69,0.0000,-1044.9,-1515.4,-743.83,-1178.1
1549.000000000,81.621,1822.3,1879.2,1059.5,264.75,2138.8,967.75,2.2765,5124.8,2738.0,3366.7,2076.0,0.0000,-6202.9,-6674.8,-1009.4,-1925.5,-1449.4,-15178.,-97.163,-18837.,-6051.1,-3924.5,-2219.3,63.629,2139.7,1950.8,1096.8,294.65,2245.0,1686.6,2.7693,6164.0,4450.3,4253.4,3658.6,0.0000,-325.14,-98.172,-67.284,-39.984,-53.285,-587.69,-0.12644,-1044.8,-1515.3,-743.80,-1178.0
1550.000000000,81.706,1823.7,1878.9,1055.0,265.13,2129.6,967.75,2.2769,5118.6,2738.0,3366.8,2076.0,0.0000,-6197.3,-6672.2,-1007.5,-1924.6,-1445.5,-15176.,-97.132,-18834.,-6050.7,-3924.1,-2218.8,59.953,2135.8,1947.5,1092.6,293.90,2235.7,1686.6,0.0000,6158.1,4449.7,4252.8,3658.0,0.0000,-324.92,-98.033,-67.154,-39.969,-53.007,-587.69,0.0000,-1044.8,-1515.3,-743.77,-1177.9
1551.000000000,81.739,1823.7,1878.8,1051.7,264.78,2121.5,967.75,2.2773,5112.5,2738.0,3366.8,2076.1,0.0000,-6192.1,-6669.9,-1005.5,-1923.6,-1441.6,-15174.,-97.101,-18832.,-6050.3,-3923.7,-2218.3,59.839,2131.7,1943.8,1088.2,293.30,2225.5,1686.6,0.0000,6152.0,4449.7,4252.8,3658.0,0.0000,-324.20,-97.797,-66.940,-39.893,-52.695,-587.69,0.0000,-1044.7,-1515.2,-743.74,-1177.8
1552.000000000,81.653,1821.6,1876.1,1048.9,264.71,2113.4,967.75,2.2778,5106.8,2738.1,3366.8,2076.2,0.0000,-6186.9,-6667.6,-1003.5,-1922.7,-1437.7,-15172.,-97.070,-18830.,-6049.9,-3923.3,-2217.8,59.657,2125.3,1937.9,1083.0,292.38,2214.1,1686.6,0.0000,6145.0,4449.7,4252.8,3658.0,0.0000,-323.10,-97.449,-66.666,-39.772,-52.354,-587.69,0.0000,-1044.6,-1515.1,-743.72,-1177.7
1553.000000000,81.652,1824.2,1878.0,1045.4,265.40,2105.2,967.75,2.2782,5101.4,2738.2,3366.8,2076.3,0.0000,-6182.1,-6665.6,-1001.6,-1921.8,-1433.9,-15171.,-97.041,-18828.,-6049.6,-3922.9,-2217.4,96.521,2216.4,2008.9,1108.1,306.39,2248.0,1686.6,47.735,6168.0,4458.8,4261.2,3667.2,0.0000,-330.47,-100.21,-67.901,-40.730,-52.970,-587.69,-2.1795,-1044.7,-1515.1,-743.73,-1177.7
1554.000000000,82.383,1840.3,1890.9,1043.0,268.16,2099.1,967.75,2.2786,5096.5,2738.2,3366.8,2076.4,0.0000,-6178.5,-6664.4,-999.86,-1921.0,-1430.1,-15169.,-97.011,-18825.,-6049.2,-3922.5,-2216.9,61.605,2194.6,2001.1,1100.4,301.62,2236.9,1686.6,0.0000,6158.8,4449.9,4252.9,3658.1,0.0000,-333.45,-100.56,-68.228,-41.070,-52.781,-587.69,0.0000,-1044.5,-1515.0,-743.66,-1177.5
1555.000000000,82.932,1854.5,1904.2,1043.1,269.39,2094.4,967.75,2.2791,5091.7,2738.2,3366.8,2076.5,0.0000,-6175.8,-6663.7,-998.12,-1920.4,-1426.3,-15167.,-96.981,-18823.,-6048.8,-3922.1,-2216.4,61.643,2196.0,2002.4,1096.6,301.72,2226.8,1686.6,0.0000,6152.5,4449.7,4252.8,3658.0,0.0000,-333.58,-100.59,-68.118,-41.095,-52.475,-587.69,0.0000,-1044.5,-1515.0,-743.63,-1177.4
1556.000000000,83.139,1860.3,1910.3,1044.2,270.82,2090.3,967.75,2.2795,5087.6,2738.3,3366.8,2076.6,0.0000,-6173.3,-6663.2,-996.42,-1919.7,-1422.7,-15165.,-96.951,-18821.,-6048.5,-3921.7,-2215.9,61.558,2193.0,1999.6,1092.1,301.26,2216.2,1686.6,0.0000,6146.0,4449.7,4252.8,3658.0,0.0000,-333.04,-100.42,-67.920,-41.038,-52.158,-587.69,0.0000,-1044.4,-1514.9,-743.60,-1177.3
1557.000000000,83.502,1861.1,1912.0,1043.1,271.53,2084.2,967.75,2.2799,5083.3,2738.4,3366.9,2076.7,0.0000,-6170.8,-6662.5,-994.72,-1919.0,-1419.0,-15163.,-96.920,-18819.,-6048.1,-3921.3,-2215.4,61.451,2189.2,1996.2,1088.0,300.70,2206.6,1686.6,0.0000,6140.2,4449.7,4252.8,3658.0,0.0000,-332.38,-100.22,-67.720,-40.967,-51.865,-587.69,0.0000,-1044.3,-1514.8,-743.58,-1177.2
1558.000000000,83.571,1860.2,1912.1,1041.3,271.34,2077.1,967.75,2.2803,5079.2,2738.4,3366.9,2076.8,0.0000,-6168.1,-6661.6,-992.99,-1918.3,-1415.3,-15161.,-96.888,-18816.,-6047.7,-3920.9,-2214.9,61.300,2183.8,1991.2,1083.5,299.92,2196.7,1686.6,0.0000,6134.1,4449.7,4252.8,3658.0,0.0000,-331.49,-99.945,-67.486,-40.866,-51.565,-587.69,0.0000,-1044.3,-1514.8,-743.55,-1177.1
1559.000000000,83.475,1857.6,1909.4,1039.3,270.75,2070.2,967.71,2.2807,5075.3,2738.5,3366.9,2076.9,0.0000,-6165.2,-6660.6,-991.24,-1917.5,-1411.6,-15159.,-96.857,-18814.,-6047.4,-3920.5,-2214.4,61.114,2177.2,1985.2,1078.7,298.99,2186.3,1686.6,0.0000,6127.9,4449.7,4252.8,3658.0,0.0000,-330.41,-99.613,-67.224,-40.743,-51.255,-587.69,0.0000,-1044.2,-1514.7,-743.52,-1177.0
1560.000000000,83.354,1853.9,1906.0,1036.4,269.87,2063.3,967.72,2.2812,5071.5,2738.5,3366.9,2077.0,0.0000,-6162.1,-6659.4,-989.51,-1916.7,-1407.8,-15157.,-96.825,-18812.,-6047.0,-3920.0,-2214.0,60.884,2168.9,1977.7,1073.4,297.84,2175.1,1686.6,0.0000,6121.1,4449.7,4252.8,3658.0,0.0000,-329.08,-99.205,-66.921,-40.589,-50.925,-587.69,0.0000,-1044.1,-1514.7,-743.49,-1177.0
1561.000000000,83.155,1849.2,1902.6,1033.0,268.99,2055.6,967.72,2.2816,5067.4,2738.6,3367.0,2077.1,0.0000,-6158.7,-6658.1,-987.75,-1915.9,-1404.0,-15156.,-96.794,-18809.,-6046.6,-3919.6,-2213.5,60.642,2160.3,1969.9,1068.0,296.64,2163.8,1686.6,0.0000,6114.3,4449.7,4252.8,3658.0,0.0000,-327.69,-98.778,-66.610,-40.428,-50.593,-587.69,0.0000,-1044.1,-1514.6,-743.46,-1176.9
1562.000000000,82.675,1845.6,1899.1,1029.1,268.22,2047.7,967.72,2.2820,5064.1,2738.7,3367.0,2077.2,0.0000,-6155.2,-6656.7,-985.97,-1915.1,-1400.1,-15154.,-96.763,-18807.,-6046.3,-3919.2,-2213.0,60.663,2202.0,1991.2,1084.3,307.12,2186.1,1686.6,0.0000,6131.9,4449.7,4263.2,3659.9,0.0000,-327.79,-99.220,-66.765,-40.506,-50.869,-587.69,0.0000,-1044.2,-1514.6,-743.48,-1176.8
1563.000000000,82.567,1842.8,1895.8,1026.3,267.74,2042.0,967.72,2.2824,5061.8,2738.7,3367.0,2077.3,0.0000,-6151.6,-6655.3,-984.20,-1914.3,-1396.3,-15152.,-96.732,-18805.,-6045.9,-3918.8,-2212.5,60.486,2154.8,1964.8,1068.9,295.94,2168.2,1686.6,36.748,6116.9,4456.3,4252.8,3661.1,0.0000,-326.69,-98.458,-66.546,-40.324,-50.586,-587.69,-1.6779,-1044.0,-1514.5,-743.40,-1176.7
1564.000000000,82.411,1839.5,1892.0,1024.1,267.04,2037.8,967.69,2.2828,5059.0,2738.7,3367.0,2077.4,0.0000,-6147.9,-6653.9,-982.42,-1913.5,-1392.6,-15150.,-96.702,-18803.,-6045.5,-3918.4,-2212.0,60.355,2150.1,1960.5,1065.5,295.28,2160.7,1686.6,0.0000,6112.4,4449.7,4252.8,3658.0,0.0000,-325.90,-98.208,-66.358,-40.237,-50.350,-587.69,0.0000,-1043.9,-1514.4,-743.38,-1176.6
1565.000000000,82.256,1838.5,1889.7,1021.9,266.92,2034.4,967.68,2.2832,5056.0,2738.8,3367.0,2077.5,0.0000,-6144.3,-6652.5,-980.66,-1912.7,-1388.8,-15148.,-96.672,-18801.,-6045.2,-3918.0,-2211.5,80.334,2228.4,2007.8,1095.4,320.69,2192.8,1686.6,56.670,6138.5,4466.3,4279.2,3674.7,0.0000,-327.49,-99.455,-66.608,-40.578,-50.535,-587.69,-2.5875,-1044.2,-1514.4,-743.48,-1176.7
1566.000000000,82.350,1840.1,1890.5,1019.3,267.09,2029.7,967.68,2.2836,5052.5,2738.8,3367.1,2077.6,0.0000,-6140.8,-6651.3,-978.94,-1911.9,-1385.2,-15146.,-96.642,-18798.,-6044.8,-3917.6,-2211.0,60.574,2157.9,1967.6,1065.1,296.28,2157.1,1686.6,0.0000,6110.2,4449.7,4252.8,3658.0,0.0000,-326.92,-98.500,-66.442,-40.382,-50.148,-587.69,0.0000,-1043.8,-1514.3,-743.32,-1176.4
1567.000000000,82.321,1839.7,1890.2,1018.0,266.78,2024.2,967.64,2.2840,5048.5,2738.8,3367.1,2077.6,0.0000,-6137.4,-6650.2,-977.22,-1911.1,-1381.5,-15144.,-96.611,-18796.,-6044.4,-3917.2,-2210.6,60.439,2153.1,1963.3,1061.2,295.59,2148.6,1686.6,0.0000,6105.1,4449.7,4252.8,3658.0,0.0000,-326.12,-98.258,-66.239,-40.293,-49.889,-587.69,0.0000,-1043.7,-1514.3,-743.29,-1176.3
1568.000000000,82.316,1838.1,1888.2,1016.6,266.71,2018.7,967.64,2.2844,5044.4,2738.9,3367.1,2077.7,0.0000,-6134.0,-6649.1,-975.50,-1910.4,-1377.8,-15142.,-96.581,-18794.,-6044.1,-3916.8,-2210.1,62.824,2152.5,1962.8,1058.4,295.47,2141.4,1686.6,0.0000,6100.7,4449.7,4252.8,3658.0,0.0000,-325.95,-98.210,-66.129,-40.282,-49.659,-587.69,0.0000,-1043.7,-1514.2,-743.26,-1176.2
1569.000000000,82.609,1835.8,1886.4,1014.1,266.48,2012.4,967.64,2.2848,5040.2,2738.9,3367.1,2077.8,0.0000,-6130.7,-6647.9,-973.81,-1909.6,-1374.2,-15140.,-96.550,-18792.,-6043.7,-3916.4,-2209.6,60.211,2145.0,1955.9,1053.4,294.41,2130.7,1686.6,0.0000,6094.2,4449.7,4252.8,3658.0,0.0000,-324.73,-97.842,-65.847,-40.141,-49.346,-587.69,0.0000,-1043.6,-1514.1,-743.23,-1176.1
1570.000000000,82.565,1831.9,1882.8,1011.6,265.72,2005.2,967.64,2.2852,5035.7,2739.0,3367.2,2077.9,0.0000,-6127.2,-6646.6,-972.11,-1908.8,-1370.5,-15139.,-96.519,-18789.,-6043.3,-3916.0,-2209.1,59.980,2136.8,1948.4,1048.1,293.26,2119.8,1686.6,0.0000,6087.6,4449.7,4252.8,3658.0,0.0000,-323.40,-97.442,-65.548,-39.987,-49.029,-587.69,0.0000,-1043.6,-1514.1,-743.20,-1176.0
1571.000000000,82.641,1826.8,1877.4,1008.5,264.96,1997.5,967.64,2.2845,5031.3,2739.0,3367.2,2077.9,0.0000,-6123.5,-6645.2,-970.37,-1908.0,-1366.8,-15137.,-96.488,-18787.,-6043.0,-3915.5,-2208.6,59.729,2127.8,1940.2,1042.7,292.01,2108.5,1686.6,0.0000,6080.8,4449.7,4252.8,3658.0,0.0000,-321.96,-97.008,-65.232,-39.819,-48.704,-587.69,0.0000,-1043.5,-1514.0,-743.17,-1175.9
1572.000000000,82.496,1820.5,1871.0,1004.8,264.00,1990.3,967.64,2.2826,5028.0,2739.1,3367.2,2078.0,0.0000,-6119.6,-6643.7,-968.62,-1907.1,-1363.1,-15135.,-96.457,-18785.,-6042.6,-3915.1,-2208.1,59.471,2118.6,1931.8,1037.3,290.74,2097.2,1686.6,0.0000,6074.0,4449.7,4252.8,3658.0,0.0000,-320.48,-96.563,-64.912,-39.647,-48.379,-587.69,0.0000,-1043.4,-1514.0,-743.15,-1175.8
1573.000000000,82.349,1813.8,1864.5,1000.8,262.99,1983.1,967.64,2.2830,5024.7,2739.2,3367.2,2078.1,0.0000,-6115.4,-6641.9,-966.85,-1906.3,-1359.3,-15133.,-96.426,-18783.,-6042.3,-3914.7,-2207.7,59.219,2109.6,1923.6,1031.9,289.49,2086.2,1686.6,0.0000,6067.4,4449.7,4252.8,3658.0,0.0000,-319.04,-96.126,-64.598,-39.479,-48.060,-587.69,0.0000,-1043.4,-1513.9,-743.12,-1175.7
1574.000000000,82.183,1807.6,1858.0,996.66,261.97,1976.0,967.64,2.2834,5021.1,2739.2,3367.3,2078.2,0.0000,-6111.1,-6640.1,-965.04,-1905.4,-1355.5,-15131.,-96.395,-18781.,-6041.9,-3914.3,-2207.2,59.020,2102.6,1917.2,1027.4,288.50,2076.7,1686.6,0.0000,6061.7,4449.7,4252.8,3658.0,0.0000,-317.88,-95.774,-64.340,-39.347,-47.779,-587.69,0.0000,-1043.3,-1513.8,-743.09,-1175.7
1575.000000000,81.953,1801.6,1851.4,992.58,261.01,1968.7,967.64,2.2838,5017.5,2739.3,3367.3,2078.3,0.0000,-6106.7,-6638.2,-963.23,-1904.5,-1351.7,-15129.,-96.364,-18778.,-6041.5,-3913.9,-2206.7,58.810,2095.1,1910.4,1022.8,287.46,2067.0,1686.6,0.0000,6055.8,4449.7,4252.8,3658.0,0.0000,-316.66,-95.402,-64.072,-39.207,-47.493,-587.69,0.0000,-1043.2,-1513.8,-743.06,-1175.6
1576.000000000,81.729,1795.7,1845.0,988.60,260.03,1961.2,967.64,2.2842,5013.6,2739.4,3367.3,2078.4,0.0000,-6102.1,-6636.3,-961.39,-1903.6,-1347.9,-15127.,-96.332,-18776.,-6041.2,-3913.5,-2206.2,58.571,2086.6,1902.6,1017.7,286.27,2056.6,1686.6,0.0000,6049.5,4449.7,4252.8,3658.0,0.0000,-315.28,-94.983,-63.774,-39.047,-47.190,-587.69,0.0000,-1043.2,-1513.7,-743.03,-1175.5
1577.000000000,81.303,1789.5,1838.7,984.46,258.93,1953.2,967.64,2.2846,5009.4,2739.4,3367.3,2078.5,0.0000,-6097.4,-6634.2,-959.53,-1902.7,-1344.1,-15125.,-96.301,-18774.,-6040.8,-3913.1,-2205.7,58.302,2077.0,1893.8,1012.2,284.94,2045.4,1686.6,0.0000,6042.7,4449.7,4252.8,3658.0,0.0000,-313.73,-94.513,-63.447,-38.868,-46.868,-587.69,0.0000,-1043.1,-1513.7,-743.00,-1175.4
1578.000000000,80.978,1782.3,1832.6,980.31,257.85,1944.7,967.64,2.2850,5004.8,2739.5,3367.3,2078.5,0.0000,-6092.5,-6632.1,-957.66,-1901.8,-1340.3,-15123.,-96.270,-18772.,-6040.4,-3912.7,-2205.2,58.070,2068.7,1886.3,1007.3,283.80,2035.2,1686.6,0.0000,6036.6,4449.7,4252.8,3658.0,0.0000,-312.39,-94.105,-63.158,-38.714,-46.572,-587.69,0.0000,-1043.1,-1513.6,-742.97,-1175.3
1579.000000000,80.798,1775.8,1826.5,975.92,256.83,1936.0,967.63,2.2853,4999.7,2739.5,3367.3,2078.6,0.0000,-6087.6,-6629.9,-955.78,-1900.8,-1336.4,-15121.,-96.239,-18769.,-6040.1,-3912.3,-2204.8,57.831,2060.2,1878.6,1002.3,282.61,2024.8,1686.6,0.0000,6030.3,4449.7,4252.8,3658.0,0.0000,-311.00,-93.682,-62.862,-38.554,-46.271,-587.69,0.0000,-1043.0,-1513.5,-742.94,-1175.2
1580.000000000,80.690,1769.1,1819.7,971.40,255.75,1927.2,967.62,2.2857,4994.5,2739.5,3367.3,2078.7,0.0000,-6082.5,-6627.6,-953.88,-1899.9,-1332.6,-15120.,-96.207,-18767.,-6039.7,-3911.8,-2204.3,57.552,2050.3,1869.5,996.67,281.24,2013.4,1686.6,0.0000,6023.5,4449.7,4252.8,3658.0,0.0000,-309.40,-93.195,-62.526,-38.368,-45.947,-587.69,0.0000,-1042.9,-1513.5,-742.91,-1175.1
1581.000000000,80.425,1761.9,1812.6,966.93,254.66,1918.0,967.62,2.2861,4989.1,2739.6,3367.4,2078.9,0.0000,-6077.4,-6625.2,-951.97,-1898.9,-1328.7,-15118.,-96.176,-18765.,-6039.3,-3911.4,-2203.8,57.337,2042.6,1862.5,992.01,280.17,2003.8,1686.6,0.0000,6017.6,4449.7,4252.8,3658.0,0.0000,-308.14,-92.811,-62.254,-38.225,-45.663,-587.69,0.0000,-1042.9,-1513.4,-742.88,-1175.0
1582.000000000,80.198,1755.2,1806.0,962.52,253.68,1908.6,967.62,2.2865,4983.7,2739.6,3367.4,2079.0,0.0000,-6072.2,-6622.9,-950.06,-1898.0,-1324.8,-15116.,-96.145,-18763.,-6039.0,-3911.0,-2203.3,57.142,2035.6,1856.2,987.66,279.20,1994.7,1686.6,0.0000,6012.1,4449.7,4252.8,3658.0,0.0000,-306.99,-92.459,-62.003,-38.094,-45.394,-587.69,0.0000,-1042.8,-1513.4,-742.86,-1174.9
1583.000000000,80.055,1748.9,1800.4,957.97,252.70,1899.8,967.62,2.2869,4978.2,2739.7,3367.4,2079.1,0.0000,-6066.9,-6620.4,-948.13,-1897.0,-1321.0,-15114.,-96.114,-18760.,-6038.6,-3910.6,-2202.8,56.917,2027.6,1848.9,982.89,278.09,1984.8,1686.6,0.0000,6006.2,4449.7,4252.8,3658.0,0.0000,-305.68,-92.058,-61.723,-37.945,-45.106,-587.69,0.0000,-1042.8,-1513.3,-742.83,-1174.8
1584.000000000,79.660,1742.3,1794.0,953.57,251.72,1891.0,967.62,2.2872,4972.9,2739.7,3367.4,2079.1,0.0000,-6061.5,-6618.0,-946.20,-1896.0,-1317.1,-15112.,-96.083,-18758.,-6038.2,-3910.2,-2202.4,56.680,2019.2,1841.2,977.92,276.91,1974.6,1686.6,0.0000,6000.0,4449.7,4252.8,3658.0,0.0000,-304.29,-91.637,-61.430,-37.787,-44.811,-587.69,0.0000,-1042.7,-1513.3,-742.80,-1174.7
1585.000000000,79.324,1735.6,1787.1,949.25,250.77,1882.2,967.62,2.2876,4967.7,2739.8,3367.5,2079.2,0.0000,-6056.1,-6615.5,-944.26,-1895.0,-1313.2,-15110.,-96.052,-18756.,-6037.9,-3909.8,-2201.9,56.455,2011.2,1833.8,973.13,275.79,1964.7,1686.6,0.0000,5994.0,4449.7,4252.8,3658.0,0.0000,-302.98,-91.235,-61.149,-37.636,-44.524,-587.69,0.0000,-1042.7,-1513.2,-742.77,-1174.6
1586.000000000,79.103,1728.9,1779.8,944.72,249.84,1873.4,967.62,2.2880,4962.6,2739.8,3367.5,2079.3,0.0000,-6050.6,-6612.9,-942.31,-1894.1,-1309.3,-15108.,-96.021,-18754.,-6037.5,-3909.4,-2201.4,56.261,2004.3,1827.6,968.82,274.83,1955.6,1686.6,0.0000,5988.6,4449.7,4252.8,3658.0,0.0000,-301.83,-90.884,-60.899,-37.507,-44.257,-587.69,0.0000,-1042.6,-1513.1,-742.74,-1174.5
1587.000000000,78.890,1722.6,1773.4,940.30,248.94,1864.5,967.59,2.2884,4957.2,2739.9,3367.5,2079.4,0.0000,-6045.0,-6610.3,-940.36,-1893.1,-1305.4,-15106.,-95.990,-18751.,-6037.2,-3909.0,-2200.9,56.059,1997.1,1821.0,964.40,273.83,1946.4,1686.6,0.0000,5983.0,4449.7,4252.8,3658.0,0.0000,-300.64,-90.520,-60.643,-37.373,-43.987,-587.69,0.0000,-1042.5,-1513.1,-742.71,-1174.4
1588.000000000,78.501,1716.4,1767.0,936.07,248.03,1855.8,967.58,2.2887,4951.8,2739.9,3367.6,2079.5,0.0000,-6039.3,-6607.7,-938.40,-1892.1,-1301.5,-15104.,-95.959,-18749.,-6036.8,-3908.5,-2200.4,55.841,1989.3,1813.9,959.73,272.75,1936.8,1686.6,0.0000,5977.2,4449.7,4252.8,3658.0,0.0000,-299.35,-90.129,-60.370,-37.227,-43.707,-587.69,0.0000,-1042.5,-1513.0,-742.68,-1174.3
1589.000000000,78.186,1710.0,1760.1,931.81,247.06,1847.3,967.59,2.2891,4946.5,2739.9,3367.6,2079.6,0.0000,-6033.6,-6605.1,-936.44,-1891.1,-1297.6,-15103.,-95.928,-18747.,-6036.4,-3908.1,-2199.9,55.616,1981.3,1806.6,954.96,271.64,1926.9,1686.6,0.0000,5971.3,4449.7,4252.8,3658.0,0.0000,-298.04,-89.728,-60.090,-37.077,-43.423,-587.69,0.0000,-1042.4,-1513.0,-742.65,-1174.2
1590.000000000,77.960,1703.7,1753.7,927.51,246.09,1838.5,967.59,2.2752,4941.2,2740.0,3367.6,2079.7,0.0000,-6027.9,-6602.4,-934.48,-1890.1,-1293.8,-15101.,-95.897,-18745.,-6036.1,-3907.7,-2199.5,55.408,1973.9,1799.9,950.46,270.60,1917.6,1686.6,0.0000,5965.6,4449.7,4252.8,3658.0,0.0000,-296.81,-89.353,-59.827,-36.939,-43.150,-587.69,0.0000,-1042.4,-1512.9,-742.62,-1174.1
1591.000000000,77.729,1697.5,1747.4,923.25,245.16,1829.6,967.56,2.2553,4935.7,2740.0,3367.6,2079.8,0.0000,-6022.1,-6599.8,-932.51,-1889.1,-1289.8,-15099.,-95.866,-18742.,-6035.7,-3907.3,-2199.0,55.185,1965.9,1792.6,945.72,269.50,1907.8,1686.6,0.0000,5959.7,4449.7,4252.8,3658.0,0.0000,-295.50,-88.953,-59.549,-36.790,-42.868,-587.69,0.0000,-1042.3,-1512.8,-742.59,-1174.0
1592.000000000,77.510,1692.9,1742.4,918.98,244.50,1821.1,967.55,2.2557,4930.6,2740.1,3367.6,2079.9,0.0000,-6016.3,-6597.2,-930.56,-1888.0,-1285.9,-15097.,-95.836,-18740.,-6035.3,-3906.9,-2198.5,56.988,1977.4,1804.4,951.92,273.61,1917.5,1686.6,0.0000,5965.8,4450.3,4255.8,3660.4,0.0000,-296.68,-89.390,-59.784,-36.969,-42.983,-587.69,0.0000,-1042.3,-1512.8,-742.58,-1174.0
1593.000000000,77.470,1691.9,1740.6,915.14,244.48,1813.6,967.55,2.2561,4925.6,2740.1,3367.6,2080.0,0.0000,-6010.8,-6594.7,-928.64,-1887.1,-1282.0,-15095.,-95.806,-18738.,-6035.0,-3906.5,-2198.0,55.330,1971.1,1797.3,945.96,270.17,1906.8,1686.6,0.0000,5959.1,4449.7,4252.8,3658.0,0.0000,-296.05,-89.113,-59.618,-36.887,-42.739,-587.69,0.0000,-1042.2,-1512.7,-742.53,-1173.9
1594.000000000,77.427,1690.1,1738.8,912.17,243.86,1806.5,967.55,2.2564,4920.7,2740.2,3367.6,2080.1,0.0000,-6005.5,-6592.4,-926.73,-1886.1,-1278.2,-15093.,-95.776,-18736.,-6034.6,-3906.1,-2197.5,55.193,1966.2,1792.9,942.11,269.47,1898.3,1686.6,0.0000,5953.9,4449.7,4252.8,3658.0,0.0000,-295.21,-88.857,-59.414,-36.795,-42.488,-587.69,0.0000,-1042.1,-1512.7,-742.50,-1173.8
1595.000000000,77.272,1686.7,1735.3,909.50,243.59,1800.0,967.55,2.2568,4916.2,2740.2,3367.6,2080.2,0.0000,-6000.2,-6590.2,-924.81,-1885.2,-1274.3,-15091.,-95.746,-18733.,-6034.3,-3905.7,-2197.1,55.024,1960.2,1787.4,937.90,268.63,1889.3,1686.6,0.0000,5948.5,4449.7,4252.8,3658.0,0.0000,-294.20,-88.549,-59.182,-36.683,-42.226,-587.69,0.0000,-1042.1,-1512.6,-742.47,-1173.7
1596.000000000,77.246,1682.3,1730.4,906.51,243.14,1793.0,967.55,2.2572,4911.7,2740.3,3367.7,2080.2,0.0000,-5994.9,-6587.9,-922.91,-1884.2,-1270.5,-15089.,-95.715,-18731.,-6033.9,-3905.2,-2196.6,54.822,1953.0,1780.8,933.28,267.62,1879.5,1686.6,0.0000,5942.6,4449.7,4252.8,3658.0,0.0000,-293.01,-88.188,-58.920,-36.548,-41.948,-587.69,0.0000,-1042.0,-1512.5,-742.45,-1173.6
1597.000000000,76.940,1677.1,1725.4,903.18,242.39,1785.6,967.55,2.2575,4906.9,2740.3,3367.7,2080.4,0.0000,-5989.5,-6585.5,-921.00,-1883.3,-1266.6,-15087.,-95.685,-18729.,-6033.5,-3904.8,-2196.1,54.621,1945.8,1774.3,928.74,266.62,1870.0,1686.6,0.0000,5936.9,4449.7,4252.8,3658.0,0.0000,-291.82,-87.829,-58.660,-36.414,-41.675,-587.69,0.0000,-1042.0,-1512.5,-742.42,-1173.5
1598.000000000,76.599,1671.7,1719.5,899.94,241.64,1778.1,967.55,2.2579,4902.4,2740.4,3367.7,2080.5,0.0000,-5984.1,-6583.1,-919.08,-1882.3,-1262.7,-15085.,-95.654,-18727.,-6033.2,-3904.4,-2195.6,54.441,1939.4,1768.4,924.42,265.72,1860.8,1686.6,0.0000,5931.3,4449.7,4252.8,3658.0,0.0000,-290.75,-87.503,-58.419,-36.294,-41.410,-587.69,0.0000,-1041.9,-1512.4,-742.39,-1173.4
1599.000000000,76.380,1666.4,1714.1,896.34,240.83,1770.2,967.55,2.2582,4897.7,2740.5,3367.8,2080.6,0.0000,-5978.5,-6580.7,-917.15,-1881.3,-1258.8,-15084.,-95.624,-18724.,-6032.8,-3904.0,-2195.2,54.231,1931.9,1761.6,919.80,264.67,1851.2,1686.6,0.0000,5925.5,4449.7,4252.8,3658.0,0.0000,-289.51,-87.129,-58.152,-36.154,-41.135,-587.69,0.0000,-1041.9,-1512.4,-742.36,-1173.3
1600.000000000,76.180,1660.6,1708.3,892.54,239.98,1762.2,967.54,2.2586,4893.1,2740.5,3367.8,2080.7,0.0000,-5972.9,-6578.3,-915.25,-1880.3,-1254.9,-15082.,-95.593,-18722.,-6032.5,-3903.6,-2194.7,54.002,1923.8,1754.2,914.94,263.54,1841.1,1686.6,0.0000,5919.4,4449.7,4252.8,3658.0,0.0000,-288.18,-86.724,-57.868,-36.001,-40.852,-587.69,0.0000,-1041.8,-1512.3,-742.33,-1173.2
1601.000000000,75.964,1656.7,1704.2,888.75,239.40,1754.2,967.54,2.2590,4888.4,2740.5,3367.8,2080.7,0.0000,-5967.4,-6575.9,-913.35,-1879.3,-1251.0,-15080.,-95.564,-18720.,-6032.1,-3903.2,-2194.2,56.805,1942.7,1769.8,927.20,270.28,1861.2,1686.6,6.3948,5932.4,4452.2,4259.6,3663.9,0.0000,-289.79,-87.314,-58.238,-36.246,-41.136,-587.69,-0.29198,-1041.8,-1512.2,-742.33,-1173.2
1602.000000000,75.959,1657.5,1703.7,885.34,239.67,1747.6,967.54,2.2597,4884.2,2740.6,3367.8,2080.8,0.0000,-5962.2,-6573.7,-911.49,-1878.4,-1247.1,-15078.,-95.535,-18717.,-6031.7,-3902.8,-2193.7,54.363,1936.6,1765.9,920.54,265.29,1851.7,1686.6,0.0000,5926.3,4450.5,4254.7,3660.0,0.0000,-289.89,-87.236,-58.224,-36.242,-40.993,-587.69,0.0000,-1041.7,-1512.2,-742.28,-1173.0
1603.000000000,75.997,1661.5,1706.6,883.04,239.91,1742.5,967.55,2.2647,4881.0,2740.6,3367.8,2080.9,0.0000,-5957.4,-6571.9,-909.68,-1877.5,-1243.3,-15076.,-95.508,-18715.,-6031.4,-3902.4,-2193.3,71.042,2006.7,1817.5,949.24,285.30,1887.3,1686.6,274.02,5955.4,4465.7,4279.6,3683.0,0.0000,-293.91,-89.003,-58.879,-36.851,-41.330,-587.69,-12.512,-1042.0,-1512.1,-742.37,-1173.3
1604.000000000,76.223,1671.1,1714.1,881.85,241.72,1739.5,967.55,2.2651,4877.7,2740.7,3367.9,2081.0,0.0000,-5953.4,-6570.5,-907.93,-1876.7,-1239.5,-15074.,-95.480,-18713.,-6031.0,-3901.9,-2192.8,55.418,1974.2,1800.2,928.37,270.27,1860.7,1686.6,0.0000,5931.8,4454.8,4261.8,3670.4,0.0000,-295.32,-88.876,-59.015,-36.945,-41.084,-587.69,0.0000,-1041.7,-1512.1,-742.25,-1173.0
1605.000000000,76.496,1679.1,1721.5,881.69,242.67,1736.9,967.55,2.2655,4874.9,2740.8,3367.9,2081.1,0.0000,-5949.9,-6569.5,-906.22,-1876.0,-1235.8,-15072.,-95.451,-18711.,-6030.7,-3901.5,-2192.3,55.452,1975.4,1801.3,926.36,270.39,1854.5,1686.6,0.0000,5927.3,4450.3,4253.6,3659.1,0.0000,-295.41,-88.907,-58.960,-36.968,-40.901,-587.69,0.0000,-1041.7,-1512.0,-742.19,-1172.7
1606.000000000,76.606,1682.5,1725.4,881.54,243.40,1734.4,967.55,2.2659,4871.5,2740.8,3367.9,2081.2,0.0000,-5946.6,-6568.6,-904.52,-1875.3,-1232.2,-15070.,-95.422,-18708.,-6030.3,-3901.1,-2191.8,55.376,1972.7,1798.8,922.98,269.98,1846.5,1686.6,0.0000,5922.5,4449.8,4252.9,3658.2,0.0000,-294.91,-88.763,-58.805,-36.917,-40.669,-587.69,0.0000,-1041.6,-1512.0,-742.15,-1172.6
1607.000000000,76.836,1682.6,1725.6,881.34,243.76,1730.5,967.55,2.2662,4868.4,2740.9,3367.9,2081.2,0.0000,-5943.2,-6567.6,-902.83,-1874.5,-1228.5,-15068.,-95.392,-18706.,-6030.0,-3900.7,-2191.4,55.219,1967.1,1793.7,918.82,269.19,1837.5,1686.6,0.0000,5917.0,4449.7,4252.8,3658.0,0.0000,-293.99,-88.490,-58.582,-36.813,-40.412,-587.69,0.0000,-1041.6,-1511.9,-742.12,-1172.5
1608.000000000,76.853,1680.3,1723.9,880.06,243.44,1725.6,967.55,2.2666,4864.6,2740.9,3368.0,2081.3,0.0000,-5939.7,-6566.5,-901.13,-1873.7,-1224.9,-15066.,-95.362,-18704.,-6029.6,-3900.3,-2190.9,55.023,1960.2,1787.3,914.30,268.22,1828.0,1686.6,0.0000,5911.2,4449.7,4252.8,3658.0,0.0000,-292.86,-88.153,-58.327,-36.682,-40.145,-587.69,0.0000,-1041.6,-1511.8,-742.09,-1172.5
1609.000000000,76.741,1676.6,1720.6,878.42,242.82,1719.7,967.53,2.2669,4861.1,2741.0,3368.0,2081.4,0.0000,-5936.1,-6565.1,-899.44,-1872.9,-1221.2,-15064.,-95.332,-18702.,-6029.3,-3899.9,-2190.4,54.815,1952.8,1780.6,909.74,267.18,1818.5,1686.6,0.0000,5905.5,4449.7,4252.8,3658.0,0.0000,-291.66,-87.797,-58.064,-36.544,-39.879,-587.69,0.0000,-1041.6,-1511.8,-742.06,-1172.4
1610.000000000,76.579,1683.2,1726.0,876.21,243.72,1713.5,967.51,2.2673,4857.4,2741.1,3368.0,2081.5,0.0000,-5932.9,-6564.2,-897.83,-1872.2,-1217.5,-15063.,-95.303,-18700.,-6028.9,-3899.5,-2189.9,180.84,2237.3,1976.0,951.98,298.64,1864.1,1686.6,15.522,5942.2,4449.7,4252.8,3658.0,0.0000,-305.40,-94.262,-59.974,-38.358,-40.361,-587.69,-0.70874,-1041.9,-1511.7,-742.03,-1172.3
1611.000000000,77.496,1714.0,1752.1,874.15,248.93,1708.3,967.51,2.2677,4853.9,2741.1,3368.0,2081.6,0.0000,-5931.8,-6564.5,-896.34,-1871.7,-1213.7,-15061.,-95.275,-18697.,-6028.5,-3899.0,-2189.5,58.486,2083.5,1899.8,932.03,284.46,1834.4,1686.6,0.0000,5914.4,4449.7,4252.8,3658.0,0.0000,-311.07,-93.665,-60.682,-38.991,-40.123,-587.69,0.0000,-1041.5,-1511.7,-742.00,-1172.2
1612.000000000,78.591,1773.8,1808.3,875.60,256.37,1706.2,967.52,2.2681,4852.4,2741.2,3368.1,2081.7,0.0000,-5934.3,-6567.3,-895.23,-1871.6,-1210.1,-15059.,-95.251,-18695.,-6028.2,-3898.6,-2189.0,2068.8,5399.3,3951.9,1067.8,362.42,2026.5,1687.0,1056.1,6047.9,4470.0,4282.6,3687.7,0.0000,-354.14,-144.06,-67.198,-44.076,-43.459,-587.69,-48.218,-1042.2,-1511.6,-742.12,-1172.5
1613.000000000,82.145,1881.1,1901.0,882.08,273.67,1714.3,967.52,2.2685,4852.9,2741.2,3368.1,2081.8,0.0000,-5942.7,-6573.8,-894.52,-1872.3,-1206.8,-15057.,-95.228,-18693.,-6027.8,-3898.2,-2188.5,156.68,2531.8,2309.6,1527.2,490.17,2412.8,1693.2,52.078,6556.3,4854.2,4636.8,4030.6,0.0000,-360.43,-110.93,-68.574,-46.143,-45.172,-587.78,-2.3778,-1049.2,-1511.6,-743.81,-1177.4
1614.000000000,85.397,1957.8,1979.3,898.79,281.91,1726.3,967.52,2.2689,4855.8,2741.3,3369.0,2082.1,0.0000,-5954.1,-6582.3,-894.00,-1873.2,-1203.7,-15055.,-95.204,-18691.,-6027.5,-3897.8,-2188.1,68.520,2441.0,2225.8,1072.3,401.27,2036.3,1686.6,0.0000,6023.5,4449.7,4272.6,3681.2,0.0000,-364.61,-109.97,-69.054,-46.106,-43.400,-587.69,0.0000,-1041.8,-1511.5,-742.01,-1172.3
1615.000000000,87.247,1999.1,2023.0,916.21,292.12,1742.5,967.52,2.2693,4858.6,2741.3,3369.2,2082.2,0.0000,-5965.8,-6590.5,-893.45,-1874.1,-1200.9,-15053.,-95.178,-18689.,-6027.2,-3897.4,-2187.6,120.50,2584.1,2236.1,1051.1,361.68,2002.0,1686.6,27.232,6009.3,4449.7,4262.1,3667.7,0.0000,-365.89,-110.45,-69.137,-45.977,-43.159,-587.69,-1.2434,-1041.6,-1511.4,-741.93,-1172.0
1616.000000000,89.313,2025.8,2052.6,927.03,297.86,1753.5,967.52,2.2697,4862.1,2741.4,3368.8,2082.2,0.0000,-5977.5,-6598.1,-892.96,-1874.8,-1198.5,-15051.,-95.151,-18687.,-6026.8,-3897.0,-2187.1,682.17,3119.4,2854.6,1277.4,516.66,2201.7,1686.6,81.635,6008.7,4640.4,4479.4,3894.3,0.0000,-373.71,-124.94,-70.092,-47.764,-44.126,-587.69,-3.7273,-1041.5,-1511.4,-742.96,-1175.2
1617.000000000,90.352,2057.0,2086.6,933.25,301.93,1760.0,967.52,2.2700,4863.1,2741.5,3369.5,2082.6,0.0000,-5989.5,-6605.7,-892.48,-1875.5,-1195.9,-15049.,-95.123,-18684.,-6026.5,-3896.6,-2186.7,70.699,2518.6,2296.6,1055.3,353.25,1990.7,1686.6,0.0000,6006.5,4449.7,4255.9,3662.8,0.0000,-376.63,-113.78,-70.531,-47.200,-43.130,-587.69,0.0000,-1041.5,-1511.3,-741.84,-1171.7
1618.000000000,91.047,2079.5,2110.8,943.60,303.81,1764.4,967.52,2.2704,4864.1,2742.4,3370.3,2082.9,0.0000,-6001.2,-6613.1,-891.98,-1876.1,-1193.1,-15047.,-95.095,-18682.,-6026.1,-3896.2,-2186.2,70.647,2516.8,2294.9,1044.5,346.56,1976.5,1686.6,0.0000,5997.7,4449.7,4252.9,3658.4,0.0000,-376.51,-113.80,-70.429,-47.126,-42.934,-587.69,0.0000,-1041.4,-1511.3,-741.80,-1171.6
1619.000000000,91.397,2092.1,2128.8,950.20,305.06,1767.0,967.52,2.2708,4863.8,2742.8,3372.3,2083.4,0.0000,-6012.4,-6619.8,-891.39,-1876.6,-1190.3,-15045.,-95.066,-18680.,-6025.8,-3895.8,-2185.7,70.440,2509.4,2288.1,1035.6,341.38,1967.8,1686.6,0.0000,5993.1,4449.7,4252.8,3658.0,0.0000,-375.57,-113.57,-70.219,-46.962,-42.757,-587.69,0.0000,-1041.3,-1511.2,-741.77,-1171.5
1620.000000000,91.596,2096.7,2139.1,954.12,305.23,1767.9,967.52,2.2711,4865.6,2744.1,3373.2,2083.1,0.0000,-6022.7,-6625.6,-890.96,-1877.0,-1187.5,-15043.,-95.037,-18678.,-6025.4,-3895.4,-2185.3,70.158,2499.3,2279.0,1031.6,339.70,1961.9,1686.6,0.0000,5989.6,4449.7,4252.8,3658.0,0.0000,-374.22,-113.20,-69.957,-46.772,-42.586,-587.69,0.0000,-1041.3,-1511.2,-741.74,-1171.4
1621.000000000,91.652,2098.8,2142.1,957.43,304.34,1766.0,967.52,2.2715,4867.2,2744.7,3371.8,2083.3,0.0000,-6031.9,-6630.7,-890.34,-1877.3,-1184.6,-15042.,-95.007,-18676.,-6025.1,-3895.0,-2184.8,69.830,2487.6,2268.3,1027.8,338.12,1955.8,1686.6,0.0000,5985.9,4449.7,4252.8,3658.0,0.0000,-372.61,-112.75,-69.658,-46.553,-42.409,-587.69,0.0000,-1041.3,-1511.1,-741.72,-1171.3
1622.000000000,91.581,2094.6,2136.2,961.43,303.01,1764.8,967.52,2.2718,4871.0,2743.8,3370.7,2083.8,0.0000,-6039.7,-6635.1,-889.61,-1877.4,-1181.6,-15040.,-94.977,-18674.,-6024.8,-3894.6,-2184.3,69.473,2474.9,2256.7,1023.8,336.42,1949.3,1686.6,0.0000,5982.1,4449.7,4252.8,3658.0,0.0000,-370.84,-112.24,-69.337,-46.315,-42.225,-587.69,0.0000,-1041.3,-1511.1,-741.69,-1171.2
1623.000000000,91.978,2092.2,2130.8,961.47,301.59,1767.3,967.52,2.2722,4878.4,2745.6,3371.1,2084.2,0.0000,-6046.3,-6639.0,-888.80,-1877.5,-1178.6,-15038.,-94.947,-18672.,-6024.5,-3894.2,-2183.8,69.107,2461.9,2244.8,1019.7,334.67,1942.8,1686.6,0.0000,5978.2,4449.7,4252.8,3658.0,0.0000,-369.00,-111.71,-69.009,-46.071,-42.039,-587.69,0.0000,-1041.2,-1511.0,-741.66,-1171.1
1624.000000000,91.248,2089.8,2127.6,959.23,300.02,1773.6,967.52,2.2725,4885.7,2746.4,3371.0,2084.7,0.0000,-6051.8,-6642.4,-887.92,-1877.6,-1175.6,-15036.,-94.917,-18670.,-6024.2,-3893.8,-2183.4,68.736,2448.7,2232.8,1015.5,332.90,1936.2,1686.6,0.0000,5974.3,4449.7,4252.8,3658.0,0.0000,-367.13,-111.17,-68.677,-45.824,-41.853,-587.69,0.0000,-1041.2,-1511.0,-741.64,-1171.1
1625.000000000,90.884,2082.5,2121.7,957.16,298.54,1777.6,967.52,2.2728,4889.8,2746.5,3370.4,2084.9,0.0000,-6056.3,-6645.3,-886.99,-1877.5,-1172.6,-15034.,-94.888,-18668.,-6024.0,-3893.4,-2182.9,68.356,2435.2,2220.5,1011.3,331.08,1929.4,1686.6,0.0000,5970.2,4449.7,4252.8,3658.0,0.0000,-365.19,-110.60,-68.336,-45.571,-41.662,-587.69,0.0000,-1041.2,-1510.9,-741.61,-1171.0
1626.000000000,90.509,2075.4,2113.6,954.93,297.10,1782.2,967.53,2.2862,4892.6,2745.8,3370.1,2085.1,0.0000,-6060.1,-6647.9,-886.00,-1877.5,-1169.5,-15032.,-94.858,-18666.,-6023.8,-3893.0,-2182.4,67.974,2421.5,2208.0,1007.0,329.25,1922.5,1686.6,0.0000,5966.1,4449.7,4252.8,3658.0,0.0000,-363.23,-110.02,-67.992,-45.316,-41.468,-587.69,0.0000,-1041.2,-1510.8,-741.59,-1170.9
1627.000000000,90.138,2066.7,2109.6,952.55,295.62,1779.9,967.53,2.9713,4894.0,2745.6,3370.1,2084.6,0.0000,-6063.6,-6650.1,-884.95,-1877.3,-1166.5,-15030.,-94.828,-18664.,-6023.5,-3892.7,-2182.0,67.588,2407.8,2195.5,1002.6,327.40,1915.5,1686.6,0.0000,5961.9,4449.7,4252.8,3658.0,0.0000,-361.23,-109.42,-67.643,-45.058,-41.271,-587.69,0.0000,-1041.1,-1510.8,-741.56,-1170.8
1628.000000000,89.760,2057.2,2102.7,950.66,294.04,1776.8,967.50,4.4673,4892.9,2743.9,3369.9,2084.5,0.0000,-6066.5,-6652.0,-883.86,-1877.2,-1163.4,-15029.,-94.798,-18662.,-6023.2,-3892.3,-2181.5,67.200,2394.0,2182.9,998.19,325.55,1908.5,1686.6,0.0000,5957.7,4449.7,4252.8,3658.0,0.0000,-359.22,-108.82,-67.294,-44.800,-41.076,-587.69,0.0000,-1041.1,-1510.7,-741.53,-1170.7
1629.000000000,89.358,2050.3,2092.6,948.08,292.41,1772.6,967.49,4.4674,4891.9,2743.7,3369.6,2084.6,0.0000,-6068.8,-6653.4,-882.73,-1876.9,-1160.3,-15027.,-94.768,-18660.,-6022.9,-3891.9,-2181.0,66.810,2380.1,2170.2,993.66,323.68,1901.1,1686.6,0.0000,5953.3,4449.7,4252.8,3658.0,0.0000,-357.18,-108.21,-66.939,-44.540,-40.873,-587.69,0.0000,-1041.1,-1510.7,-741.51,-1170.6
1630.000000000,88.473,2040.3,2082.8,944.58,290.79,1767.2,967.49,4.4675,4889.2,2743.7,3369.6,2084.8,0.0000,-6070.5,-6654.4,-881.55,-1876.6,-1157.2,-15025.,-94.739,-18658.,-6022.6,-3891.5,-2180.6,66.416,2366.0,2157.4,989.03,321.79,1893.5,1686.6,0.0000,5948.8,4449.7,4252.8,3658.0,0.0000,-355.11,-107.59,-66.579,-44.277,-40.665,-587.69,0.0000,-1041.1,-1510.6,-741.48,-1170.5
1631.000000000,88.043,2029.4,2072.4,940.97,289.18,1761.8,967.48,4.1634,4886.1,2743.8,3369.6,2084.8,0.0000,-6071.6,-6655.0,-880.34,-1876.3,-1154.1,-15023.,-94.709,-18656.,-6022.3,-3891.1,-2180.1,66.028,2352.2,2144.8,984.45,319.93,1886.0,1686.6,0.0000,5944.3,4449.7,4252.8,3658.0,0.0000,-353.07,-106.97,-66.224,-44.019,-40.458,-587.69,0.0000,-1041.0,-1510.6,-741.45,-1170.4
1632.000000000,87.654,2018.6,2061.3,938.77,287.51,1756.7,967.48,3.8981,4883.0,2743.8,3369.6,2084.8,0.0000,-6072.2,-6655.3,-879.09,-1875.9,-1151.0,-15021.,-94.679,-18654.,-6022.0,-3890.7,-2179.6,65.658,2339.0,2132.8,980.04,318.16,1878.7,1686.6,0.0000,5939.9,4449.7,4252.8,3658.0,0.0000,-351.11,-106.38,-65.883,-43.772,-40.257,-587.69,0.0000,-1041.0,-1510.5,-741.42,-1170.3
1633.000000000,87.274,2008.3,2049.8,935.68,285.92,1752.2,967.48,5.7956,4880.2,2743.9,3369.6,2085.0,0.0000,-6072.3,-6655.2,-877.80,-1875.5,-1147.9,-15019.,-94.650,-18653.,-6021.7,-3890.3,-2179.2,65.289,2325.9,2120.8,975.59,316.39,1871.3,1686.6,0.0000,5935.5,4449.7,4252.8,3658.0,0.0000,-349.15,-105.78,-65.541,-43.526,-40.054,-587.69,0.0000,-1041.0,-1510.5,-741.40,-1170.3
1634.000000000,86.970,1998.8,2038.9,932.82,284.38,1747.1,967.48,5.8586,4877.9,2743.9,3369.5,2085.1,0.0000,-6072.0,-6654.7,-876.49,-1875.0,-1144.9,-15017.,-94.620,-18651.,-6021.3,-3889.9,-2178.7,64.930,2313.1,2109.2,971.23,314.66,1864.1,1686.6,0.0000,5931.1,4449.7,4252.8,3658.0,0.0000,-347.23,-105.19,-65.208,-43.287,-39.853,-587.69,0.0000,-1041.0,-1510.4,-741.37,-1170.2
1635.000000000,86.711,1987.7,2029.5,930.62,282.86,1743.1,967.45,5.5227,4875.3,2744.0,3369.5,2085.3,0.0000,-6071.2,-6654.1,-875.15,-1874.5,-1141.8,-15016.,-94.590,-18649.,-6021.0,-3889.4,-2178.2,64.571,2300.3,2097.5,966.82,312.94,1856.6,1686.6,0.0000,5926.7,4449.7,4252.8,3658.0,0.0000,-345.30,-104.60,-64.872,-43.047,-39.650,-587.69,0.0000,-1041.0,-1510.3,-741.34,-1170.1
1636.000000000,86.348,1977.0,2020.8,927.09,281.37,1738.1,967.45,5.1659,4871.6,2744.0,3369.4,2085.3,0.0000,-6070.1,-6653.1,-873.79,-1873.9,-1138.7,-15014.,-94.561,-18647.,-6020.7,-3889.0,-2177.8,64.216,2287.7,2086.0,962.54,311.24,1849.5,1686.6,0.0000,5922.5,4449.7,4252.8,3658.0,0.0000,-343.38,-104.02,-64.544,-42.810,-39.453,-587.69,0.0000,-1040.9,-1510.3,-741.31,-1170.0
1637.000000000,85.998,1967.9,2018.2,924.30,279.91,1732.4,967.45,5.4239,4867.9,2744.2,3369.3,2085.4,0.0000,-6069.0,-6652.0,-872.41,-1873.3,-1135.6,-15012.,-94.531,-18645.,-6020.3,-3888.6,-2177.3,63.882,2275.8,2075.1,958.38,309.63,1842.5,1686.6,0.0000,5918.2,4449.7,4252.8,3658.0,0.0000,-341.58,-103.46,-64.230,-42.588,-39.258,-587.69,0.0000,-1040.9,-1510.2,-741.28,-1169.9
1638.000000000,85.659,1959.2,2008.3,920.53,278.50,1726.7,967.45,5.5395,4864.5,2744.2,3369.2,2085.3,0.0000,-6067.6,-6650.6,-871.01,-1872.7,-1132.5,-15010.,-94.502,-18643.,-6020.0,-3888.2,-2176.8,63.545,2263.8,2064.2,954.15,308.02,1835.3,1686.6,0.0000,5913.9,4449.7,4252.8,3658.0,0.0000,-339.75,-102.90,-63.912,-42.364,-39.060,-587.69,0.0000,-1040.9,-1510.2,-741.25,-1169.8
1639.000000000,85.392,1951.3,2001.0,916.69,277.43,1720.7,967.44,5.5487,4861.9,2744.5,3369.2,2085.4,0.0000,-6066.2,-6649.2,-869.61,-1872.1,-1129.4,-15008.,-94.473,-18641.,-6019.7,-3887.8,-2176.4,84.443,2298.2,2099.1,966.71,319.94,1843.0,1686.6,0.0000,5914.6,4449.7,4252.8,3658.0,0.0000,-340.52,-103.76,-64.013,-42.526,-39.073,-587.69,0.0000,-1040.9,-1510.1,-741.22,-1169.7
1640.000000000,85.335,1947.1,1998.3,915.05,277.02,1714.9,967.42,5.2537,4859.1,2744.6,3369.4,2085.5,0.0000,-6065.0,-6647.8,-868.22,-1871.5,-1126.3,-15006.,-94.444,-18639.,-6019.3,-3887.4,-2175.9,63.523,2263.0,2063.5,952.34,307.88,1830.9,1686.6,0.0000,5911.2,4449.7,4252.8,3658.0,0.0000,-339.57,-102.83,-63.832,-42.349,-38.883,-587.69,0.0000,-1040.8,-1510.1,-741.19,-1169.6
1641.000000000,85.227,1941.9,1997.3,912.55,276.11,1709.8,967.42,4.7312,4855.9,2744.6,3369.4,2085.7,0.0000,-6063.9,-6646.5,-866.82,-1871.0,-1123.3,-15005.,-94.415,-18637.,-6019.0,-3887.0,-2175.5,63.254,2253.4,2054.7,948.46,306.58,1823.8,1686.6,0.0000,5907.0,4449.7,4252.8,3658.0,0.0000,-338.10,-102.38,-63.560,-42.169,-38.688,-587.69,0.0000,-1040.8,-1510.0,-741.16,-1169.5
1642.000000000,85.016,1934.7,1991.5,910.14,275.39,1705.3,967.39,5.3449,4852.8,2744.7,3369.4,2085.7,0.0000,-6062.5,-6645.0,-865.41,-1870.3,-1120.2,-15003.,-94.386,-18635.,-6018.7,-3886.6,-2175.0,62.949,2242.5,2044.8,944.23,305.11,1816.2,1686.6,0.0000,5902.5,4449.7,4252.8,3658.0,0.0000,-336.43,-101.87,-63.259,-41.966,-38.482,-587.69,0.0000,-1040.8,-1509.9,-741.14,-1169.4
1643.000000000,84.825,1926.4,1984.0,907.23,274.40,1700.1,967.39,6.2399,4849.9,2744.8,3369.4,2085.7,0.0000,-6060.9,-6643.4,-863.98,-1869.7,-1117.2,-15001.,-94.357,-18633.,-6018.3,-3886.2,-2174.5,62.654,2232.0,2035.2,940.17,303.69,1809.0,1686.6,0.0000,5898.2,4449.7,4252.8,3658.0,0.0000,-334.81,-101.37,-62.969,-41.769,-38.284,-587.69,0.0000,-1040.8,-1509.9,-741.11,-1169.3
1644.000000000,84.440,1917.8,1975.3,903.80,273.23,1694.2,967.39,6.2400,4846.4,2745.0,3369.4,2085.7,0.0000,-6059.0,-6641.6,-862.54,-1869.0,-1114.1,-14999.,-94.327,-18631.,-6018.0,-3885.8,-2174.1,62.367,2221.8,2025.9,936.23,302.30,1802.0,1686.6,0.0000,5894.0,4449.7,4252.8,3658.0,0.0000,-333.22,-100.88,-62.687,-41.578,-38.092,-587.69,0.0000,-1040.8,-1509.8,-741.08,-1169.3
1645.000000000,83.944,1909.0,1966.6,900.55,272.02,1688.6,967.39,5.9477,4843.0,2745.2,3369.3,2085.8,0.0000,-6056.7,-6639.6,-861.08,-1868.3,-1111.1,-14997.,-94.298,-18629.,-6017.7,-3885.4,-2173.6,62.074,2211.3,2016.4,932.24,300.89,1795.0,1686.6,0.0000,5889.7,4449.7,4252.8,3658.0,0.0000,-331.60,-100.38,-62.400,-41.382,-37.897,-587.69,0.0000,-1040.7,-1509.8,-741.05,-1169.2
1646.000000000,83.638,1900.0,1958.0,897.14,270.79,1683.2,967.39,5.3118,4839.8,2745.3,3369.3,2085.9,0.0000,-6054.2,-6637.6,-859.60,-1867.6,-1108.0,-14995.,-94.269,-18627.,-6017.3,-3885.0,-2173.2,61.777,2200.8,2006.7,928.20,299.46,1787.8,1686.6,0.0000,5885.4,4449.7,4252.8,3658.0,0.0000,-329.96,-99.875,-62.109,-41.185,-37.702,-587.69,0.0000,-1040.7,-1509.7,-741.02,-1169.1
1647.000000000,83.187,1891.6,1949.5,893.66,269.61,1678.1,967.39,5.3928,4836.9,2745.3,3369.3,2086.0,0.0000,-6051.4,-6635.5,-858.11,-1866.8,-1104.8,-14994.,-94.239,-18625.,-6017.0,-3884.5,-2172.7,61.545,2192.5,1999.2,924.63,298.33,1781.2,1686.6,0.0000,5881.4,4449.7,4252.8,3658.0,0.0000,-328.66,-99.473,-61.868,-41.030,-37.517,-587.69,0.0000,-1040.7,-1509.7,-740.99,-1169.0
1648.000000000,82.816,1884.0,1941.4,890.17,268.58,1672.0,967.39,6.9111,4834.5,2744.9,3369.3,2086.0,0.0000,-6048.3,-6633.3,-856.62,-1866.1,-1101.7,-14992.,-94.210,-18623.,-6016.7,-3884.1,-2172.2,61.292,2183.5,1991.0,921.17,297.11,1775.1,1686.6,0.0000,5877.8,4449.7,4252.8,3658.0,0.0000,-327.25,-99.036,-61.619,-40.861,-37.344,-587.69,0.0000,-1040.7,-1509.6,-740.96,-1168.9
1649.000000000,82.739,1877.6,1934.5,886.87,267.69,1666.0,967.39,6.9112,4832.2,2744.8,3369.3,2086.1,0.0000,-6045.2,-6631.1,-855.12,-1865.3,-1098.5,-14990.,-94.182,-18621.,-6016.3,-3883.7,-2171.8,66.554,2183.4,1990.9,921.97,297.08,1778.6,1686.6,0.0000,5878.6,4449.7,4256.5,3658.1,0.0000,-327.16,-99.004,-61.589,-40.859,-37.289,-587.69,0.0000,-1040.7,-1509.5,-740.95,-1168.8
1650.000000000,82.592,1877.0,1932.2,883.63,267.75,1661.0,967.39,6.5027,4829.2,2744.5,3369.3,2086.2,0.0000,-6042.3,-6629.2,-853.66,-1864.6,-1095.4,-14988.,-94.154,-18619.,-6016.0,-3883.3,-2171.3,94.415,2247.4,2034.6,942.61,303.90,1800.3,1686.6,4.3073,5893.5,4453.1,4259.1,3660.0,0.0000,-330.69,-100.52,-62.101,-41.322,-37.457,-587.69,-0.19667,-1040.8,-1509.5,-740.93,-1168.7
1651.000000000,82.817,1883.2,1936.2,880.98,268.68,1657.6,967.39,6.8500,4826.6,2744.6,3369.3,2086.3,0.0000,-6040.0,-6627.8,-852.23,-1863.9,-1092.2,-14986.,-94.126,-18617.,-6015.6,-3882.9,-2170.9,62.060,2210.8,2015.9,924.87,300.70,1776.0,1686.6,0.0000,5878.2,4449.7,4252.8,3658.0,0.0000,-331.16,-100.21,-62.122,-41.373,-37.243,-587.69,0.0000,-1040.6,-1509.4,-740.87,-1168.6
1652.000000000,82.814,1886.6,1939.2,879.63,268.82,1654.3,967.39,6.6715,4824.7,2744.7,3369.3,2086.3,0.0000,-6038.1,-6626.6,-850.83,-1863.3,-1089.1,-14985.,-94.098,-18615.,-6015.3,-3882.5,-2170.4,61.948,2206.9,2012.3,922.07,300.13,1770.0,1686.6,0.0000,5874.5,4449.7,4252.8,3658.0,0.0000,-330.51,-100.01,-61.969,-41.298,-37.072,-587.69,0.0000,-1040.6,-1509.4,-740.84,-1168.5
1653.000000000,82.819,1885.3,1937.9,878.57,269.14,1651.6,967.39,5.9863,4821.8,2744.7,3369.4,2086.6,0.0000,-6036.1,-6625.4,-849.42,-1862.7,-1086.1,-14983.,-94.069,-18613.,-6014.9,-3882.1,-2170.0,61.765,2200.4,2006.4,918.81,299.24,1763.6,1686.6,0.0000,5870.7,4449.7,4252.8,3658.0,0.0000,-329.48,-99.693,-61.763,-41.177,-36.893,-587.69,0.0000,-1040.6,-1509.3,-740.81,-1168.4
1654.000000000,82.756,1881.3,1934.3,876.92,268.93,1647.8,967.39,5.9864,4819.0,2744.7,3369.4,2086.9,0.0000,-6034.0,-6624.1,-848.01,-1862.1,-1083.1,-14981.,-94.041,-18611.,-6014.6,-3881.7,-2169.5,61.547,2192.6,1999.3,915.32,298.18,1757.0,1686.6,0.0000,5866.7,4449.7,4252.8,3658.0,0.0000,-328.26,-99.321,-61.532,-41.031,-36.711,-587.69,0.0000,-1040.5,-1509.3,-740.78,-1168.3
1655.000000000,82.614,1876.2,1929.6,874.64,268.21,1643.0,967.40,5.9866,4816.0,2744.8,3369.4,2086.8,0.0000,-6031.6,-6622.6,-846.58,-1861.4,-1080.1,-14979.,-94.012,-18609.,-6014.2,-3881.3,-2169.0,61.313,2184.2,1991.7,911.78,297.04,1750.4,1686.6,0.0000,5862.8,4449.7,4252.8,3658.0,0.0000,-326.95,-98.921,-61.290,-40.875,-36.530,-587.69,0.0000,-1040.5,-1509.2,-740.75,-1168.2
1656.000000000,82.599,1871.3,1923.9,872.43,267.35,1638.2,967.40,5.3773,4812.8,2744.8,3369.5,2086.8,0.0000,-6029.0,-6621.0,-845.14,-1860.7,-1077.0,-14977.,-93.983,-18607.,-6013.9,-3880.9,-2168.6,61.134,2177.9,1985.8,908.94,296.17,1745.1,1686.6,0.0000,5859.6,4449.7,4252.8,3658.0,0.0000,-325.93,-98.611,-61.100,-40.756,-36.376,-587.69,0.0000,-1040.5,-1509.1,-740.72,-1168.2
1657.000000000,82.402,1866.2,1918.6,869.96,266.53,1633.7,967.40,5.0583,4809.5,2744.9,3369.6,2087.0,0.0000,-6026.3,-6619.4,-843.68,-1859.9,-1073.9,-14976.,-93.954,-18605.,-6013.5,-3880.5,-2168.1,60.953,2171.4,1980.0,907.15,295.31,1742.4,1686.6,0.0000,5858.0,4450.0,4253.8,3659.2,0.0000,-324.91,-98.297,-60.943,-40.635,-36.282,-587.69,0.0000,-1040.5,-1509.1,-740.70,-1168.1
1658.000000000,82.206,1861.7,1914.5,867.39,265.84,1628.7,967.40,5.2685,4806.3,2744.9,3369.7,2087.2,0.0000,-6023.5,-6617.8,-842.25,-1859.2,-1070.8,-14974.,-93.926,-18603.,-6013.2,-3880.1,-2167.7,60.992,2213.2,1984.5,923.20,295.50,1745.3,1686.6,0.0000,5862.3,4449.7,4252.8,3658.0,0.0000,-325.11,-98.407,-60.964,-40.661,-36.257,-587.69,0.0000,-1040.5,-1509.0,-740.66,-1168.0
1659.000000000,82.112,1859.4,1912.2,865.18,265.54,1624.8,967.40,6.6595,4803.4,2745.0,3369.7,2087.3,0.0000,-6020.8,-6616.2,-840.83,-1858.5,-1067.7,-14972.,-93.898,-18601.,-6012.8,-3879.7,-2167.2,60.891,2169.2,1978.0,905.86,295.01,1739.8,1686.6,0.0000,5856.4,4449.7,4252.8,3658.0,0.0000,-324.45,-98.153,-60.859,-40.594,-36.149,-587.69,0.0000,-1040.4,-1509.0,-740.63,-1167.9
1660.000000000,82.013,1858.1,1908.8,863.63,265.02,1620.8,967.40,6.6619,4800.6,2745.0,3369.7,2087.3,0.0000,-6018.0,-6614.7,-839.40,-1857.8,-1064.6,-14970.,-93.870,-18599.,-6012.5,-3879.3,-2166.7,60.722,2163.2,1972.5,903.01,294.18,1734.3,1686.6,0.0000,5853.1,4449.7,4252.8,3658.0,0.0000,-323.48,-97.858,-60.674,-40.481,-35.992,-587.69,0.0000,-1040.4,-1508.9,-740.60,-1167.8
1661.000000000,81.874,1855.3,1904.0,861.96,264.50,1616.9,967.40,6.6633,4798.3,2745.1,3369.7,2087.3,0.0000,-6015.1,-6613.1,-837.96,-1857.1,-1061.5,-14968.,-93.841,-18597.,-6012.1,-3878.9,-2166.3,60.477,2154.5,1964.5,899.58,293.00,1728.1,1686.6,0.0000,5849.4,4449.7,4252.8,3658.0,0.0000,-322.11,-97.440,-60.430,-40.318,-35.821,-587.69,0.0000,-1040.4,-1508.9,-740.57,-1167.7
1662.000000000,81.725,1849.7,1898.2,859.87,263.74,1614.1,967.40,6.3687,4796.4,2745.4,3369.7,2087.3,0.0000,-6012.1,-6611.4,-836.51,-1856.3,-1058.4,-14967.,-93.813,-18595.,-6011.8,-3878.5,-2165.8,60.218,2145.2,1956.1,895.89,291.75,1721.5,1686.6,0.0000,5845.4,4449.7,4252.8,3658.0,0.0000,-320.67,-96.999,-60.172,-40.146,-35.640,-587.69,0.0000,-1040.4,-1508.8,-740.55,-1167.6
1663.000000000,81.514,1843.0,1891.8,857.35,262.79,1610.8,967.40,6.0485,4794.1,2745.5,3369.8,2087.3,0.0000,-6008.8,-6609.7,-835.05,-1855.5,-1055.3,-14965.,-93.784,-18593.,-6011.5,-3878.1,-2165.3,59.951,2135.7,1947.4,892.11,290.46,1714.7,1686.6,0.0000,5841.3,4449.7,4252.8,3658.0,0.0000,-319.17,-96.543,-59.906,-39.968,-35.456,-587.69,0.0000,-1040.3,-1508.7,-740.52,-1167.5
1664.000000000,81.273,1836.1,1884.8,854.75,261.73,1606.6,967.40,5.1824,4792.7,2745.6,3369.9,2087.3,0.0000,-6005.3,-6607.8,-833.58,-1854.7,-1052.2,-14963.,-93.755,-18591.,-6011.1,-3877.7,-2164.9,59.681,2126.1,1938.7,888.30,289.15,1707.8,1686.6,0.0000,5837.2,4449.7,4252.8,3658.0,0.0000,-317.66,-96.081,-59.637,-39.787,-35.271,-587.69,0.0000,-1040.3,-1508.7,-740.49,-1167.4
1665.000000000,81.023,1828.8,1877.7,852.08,260.62,1602.1,967.37,5.1195,4790.0,2745.6,3369.8,2087.4,0.0000,-6001.7,-6605.9,-832.09,-1853.9,-1049.1,-14961.,-93.726,-18589.,-6010.8,-3877.3,-2164.4,59.414,2116.6,1930.0,884.50,287.86,1701.0,1686.6,0.0000,5833.1,4449.7,4252.8,3658.0,0.0000,-316.16,-95.623,-59.370,-39.609,-35.086,-587.69,0.0000,-1040.3,-1508.6,-740.46,-1167.3
1666.000000000,80.760,1830.1,1878.1,849.26,260.90,1597.1,967.37,5.1197,4787.2,2745.7,3369.9,2087.3,0.0000,-5998.5,-6604.2,-830.68,-1853.2,-1046.0,-14959.,-93.699,-18587.,-6010.4,-3876.9,-2164.0,101.15,2299.1,2011.7,916.57,299.58,1730.5,1686.6,0.0000,5853.4,4449.7,4254.6,3658.1,0.0000,-325.69,-98.969,-60.780,-40.808,-35.511,-587.69,0.0000,-1040.4,-1508.6,-740.44,-1167.2
1667.000000000,81.402,1850.0,1894.0,847.03,264.28,1593.5,967.37,5.1199,4784.6,2745.8,3369.9,2087.4,0.0000,-5996.8,-6603.6,-829.35,-1852.6,-1042.8,-14958.,-93.672,-18585.,-6010.1,-3876.5,-2163.5,61.859,2203.7,2009.4,902.80,299.39,1720.1,1686.6,0.0000,5844.2,4449.7,4252.8,3658.0,0.0000,-329.06,-99.531,-61.215,-41.239,-35.412,-587.69,0.0000,-1040.3,-1508.5,-740.40,-1167.2
1668.000000000,82.018,1867.0,1910.4,847.63,265.52,1590.8,967.37,5.1217,4783.0,2746.1,3369.9,2087.4,0.0000,-5996.1,-6603.7,-828.09,-1852.2,-1039.7,-14956.,-93.644,-18583.,-6009.8,-3876.1,-2163.0,61.899,2205.1,2010.7,900.57,299.54,1714.5,1686.6,0.0000,5840.8,4449.7,4252.8,3658.0,0.0000,-329.23,-99.588,-61.168,-41.266,-35.254,-587.69,0.0000,-1040.2,-1508.5,-740.37,-1167.1
1669.000000000,82.252,1873.7,1917.3,848.87,267.21,1588.9,967.37,5.1114,4780.6,2746.4,3369.9,2087.3,0.0000,-5995.6,-6603.9,-826.83,-1851.7,-1036.7,-14954.,-93.616,-18581.,-6009.4,-3875.7,-2162.6,61.795,2201.4,2007.3,897.79,299.02,1708.6,1686.6,0.0000,5837.3,4449.7,4252.8,3658.0,0.0000,-328.63,-99.416,-61.021,-41.197,-35.090,-587.69,0.0000,-1040.2,-1508.4,-740.34,-1167.0
1670.000000000,82.652,1874.4,1918.2,849.39,268.22,1586.7,967.37,4.9653,4778.8,2746.2,3370.0,2087.4,0.0000,-5994.9,-6603.8,-825.55,-1851.2,-1033.7,-14952.,-93.588,-18579.,-6009.1,-3875.3,-2162.1,61.623,2195.3,2001.7,894.69,298.18,1702.5,1686.6,0.0000,5833.6,4449.7,4252.8,3658.0,0.0000,-327.68,-99.132,-60.827,-41.082,-34.922,-587.69,0.0000,-1040.2,-1508.3,-740.31,-1166.9
1671.000000000,82.515,1872.0,1917.2,847.90,267.96,1583.8,967.37,4.4781,4776.9,2746.1,3370.1,2087.5,0.0000,-5994.0,-6603.5,-824.25,-1850.7,-1030.7,-14950.,-93.559,-18577.,-6008.8,-3874.9,-2161.6,61.410,2187.7,1994.8,891.34,297.14,1696.2,1686.6,0.0000,5829.8,4449.7,4252.8,3658.0,0.0000,-326.50,-98.779,-60.603,-40.940,-34.751,-587.69,0.0000,-1040.2,-1508.3,-740.28,-1166.8
1672.000000000,82.376,1868.3,1913.0,846.53,267.23,1580.5,967.37,4.4784,4774.7,2746.0,3370.1,2087.6,0.0000,-5992.7,-6603.0,-822.93,-1850.1,-1027.7,-14949.,-93.530,-18575.,-6008.4,-3874.5,-2161.2,61.173,2179.3,1987.1,887.86,295.99,1689.8,1686.6,0.0000,5826.0,4449.7,4252.8,3658.0,0.0000,-325.20,-98.389,-60.364,-40.782,-34.579,-587.69,0.0000,-1040.1,-1508.2,-740.25,-1166.7
1673.000000000,82.180,1864.1,1909.5,845.31,266.45,1576.7,967.37,4.4786,4772.7,2746.1,3370.2,2087.8,0.0000,-5991.2,-6602.3,-821.58,-1849.5,-1024.7,-14947.,-93.502,-18573.,-6008.1,-3874.1,-2160.7,61.082,2176.0,1984.2,886.17,295.55,1686.5,1686.6,0.0000,5823.9,4449.7,4252.8,3658.0,0.0000,-324.67,-98.232,-60.257,-40.722,-34.470,-587.69,0.0000,-1040.1,-1508.2,-740.23,-1166.6
1674.000000000,82.025,1860.3,1907.3,843.23,265.86,1572.7,967.37,4.4788,4770.5,2746.0,3370.2,2087.9,0.0000,-5989.5,-6601.5,-820.22,-1848.8,-1021.6,-14945.,-93.473,-18571.,-6007.8,-3873.7,-2160.3,60.932,2170.7,1979.3,883.47,294.81,1681.1,1686.6,0.0000,5820.7,4449.7,4252.8,3658.0,0.0000,-323.82,-97.978,-60.087,-40.621,-34.321,-587.69,0.0000,-1040.1,-1508.1,-740.20,-1166.5
1675.000000000,81.863,1858.8,1906.1,841.10,265.19,1568.4,967.36,4.4790,4768.7,2745.8,3370.2,2087.9,0.0000,-5987.9,-6600.6,-818.89,-1848.2,-1018.5,-14943.,-93.445,-18569.,-6007.5,-3873.3,-2159.8,99.413,2170.9,1979.5,882.15,294.82,1677.6,1686.6,0.0000,5818.6,4449.7,4252.8,3658.0,0.0000,-323.81,-97.976,-60.044,-40.626,-34.209,-587.69,0.0000,-1040.1,-1508.1,-740.17,-1166.4
1676.000000000,81.745,1857.3,1904.0,840.16,264.91,1563.7,967.35,4.4810,4766.2,2745.7,3370.2,2087.9,0.0000,-5986.2,-6599.8,-817.55,-1847.5,-1015.4,-14941.,-93.417,-18567.,-6007.1,-3872.9,-2159.3,60.890,2169.2,1977.9,881.06,294.58,1675.4,1686.6,0.0000,5817.2,4449.7,4252.8,3658.0,0.0000,-323.50,-97.883,-59.978,-40.593,-34.125,-587.69,0.0000,-1040.1,-1508.0,-740.14,-1166.3
1677.000000000,81.434,1855.1,1901.0,838.87,264.46,1559.2,967.35,4.4841,4764.1,2745.6,3370.2,2088.1,0.0000,-5984.3,-6598.9,-816.20,-1846.9,-1012.4,-14940.,-93.389,-18565.,-6006.8,-3872.5,-2158.9,60.651,2160.6,1970.1,877.69,293.42,1669.3,1686.6,0.0000,5813.6,4449.7,4252.8,3658.0,0.0000,-322.17,-97.483,-59.740,-40.434,-33.961,-587.69,0.0000,-1040.0,-1507.9,-740.11,-1166.2
1678.000000000,81.278,1851.6,1896.7,837.08,263.75,1555.3,967.35,4.5111,4762.6,2745.7,3370.2,2088.2,0.0000,-5982.2,-6597.9,-814.84,-1846.2,-1009.3,-14938.,-93.361,-18563.,-6006.4,-3872.1,-2158.4,60.399,2151.7,1962.0,874.28,292.21,1663.3,1686.6,0.0000,5810.0,4449.7,4252.8,3658.0,0.0000,-320.78,-97.062,-59.495,-40.266,-33.797,-587.69,0.0000,-1040.0,-1507.9,-740.08,-1166.2
1679.000000000,81.108,1845.8,1891.6,834.96,262.99,1552.2,967.20,4.5113,4761.2,2745.9,3370.2,2088.3,0.0000,-5979.8,-6596.8,-813.46,-1845.5,-1006.2,-14936.,-93.332,-18561.,-6006.1,-3871.7,-2158.0,60.135,2142.3,1953.4,870.69,290.93,1656.9,1686.6,0.0000,5806.2,4449.7,4252.8,3658.0,0.0000,-319.32,-96.620,-59.237,-40.090,-33.627,-587.69,0.0000,-1040.0,-1507.8,-740.05,-1166.1
1680.000000000,80.900,1839.1,1885.3,832.46,262.00,1548.6,967.20,4.5116,4759.3,2746.1,3370.3,2088.4,0.0000,-5977.2,-6595.6,-812.06,-1844.8,-1003.2,-14934.,-93.304,-18559.,-6005.7,-3871.3,-2157.5,59.874,2133.0,1944.9,867.14,289.68,1650.7,1686.6,0.0000,5802.4,4449.7,4252.8,3658.0,0.0000,-317.88,-96.181,-58.982,-39.916,-33.459,-587.69,0.0000,-1040.0,-1507.8,-740.02,-1166.0
1681.000000000,80.643,1832.7,1879.1,830.13,260.95,1545.5,967.20,4.5118,4757.2,2746.2,3370.2,2088.5,0.0000,-5974.3,-6594.2,-810.64,-1844.1,-1000.1,-14932.,-93.275,-18557.,-6005.4,-3870.9,-2157.0,59.634,2124.4,1937.1,864.00,288.52,1645.2,1686.6,0.0000,5799.2,4449.7,4252.8,3658.0,0.0000,-316.54,-95.775,-58.752,-39.756,-33.309,-587.69,0.0000,-1040.0,-1507.7,-739.99,-1165.9
1682.000000000,80.395,1849.2,1894.1,827.42,263.70,1541.4,967.20,4.5120,4754.8,2746.2,3370.2,2088.6,0.0000,-5972.9,-6593.8,-809.40,-1843.5,-997.00,-14931.,-93.249,-18555.,-6005.0,-3870.5,-2156.6,518.74,2636.6,2224.6,898.47,315.64,1663.9,1686.6,0.0000,5808.9,4450.0,4252.8,3658.6,0.0000,-343.97,-106.55,-62.329,-43.162,-33.623,-587.69,0.0000,-1039.9,-1507.7,-739.97,-1165.8
1683.000000000,82.620,1912.2,1947.0,825.71,274.01,1537.9,967.20,4.5024,4752.3,2746.4,3370.3,2088.7,0.0000,-5975.6,-6596.0,-808.31,-1843.5,-993.94,-14929.,-93.223,-18553.,-6004.7,-3870.1,-2156.1,66.302,2362.0,2153.7,898.71,321.36,1660.1,1686.6,0.0000,5806.9,4449.7,4252.8,3658.0,0.0000,-351.92,-106.52,-63.342,-44.211,-33.511,-587.69,0.0000,-1039.9,-1507.6,-739.94,-1165.7
1684.000000000,84.366,1961.5,1996.1,830.28,277.76,1534.9,967.20,3.8970,4750.1,2746.6,3370.4,2088.8,0.0000,-5980.6,-6599.9,-807.40,-1843.7,-990.91,-14927.,-93.196,-18551.,-6004.3,-3869.7,-2155.7,66.470,2367.9,2159.2,898.07,320.99,1656.6,1686.6,0.0000,5804.7,4449.7,4252.8,3658.0,0.0000,-352.84,-106.83,-63.405,-44.316,-33.399,-587.69,0.0000,-1039.9,-1507.6,-739.91,-1165.6
1685.000000000,85.214,1982.4,2018.5,835.63,283.00,1533.8,967.16,3.8968,4747.6,2746.7,3370.4,2088.9,0.0000,-5985.7,-6603.6,-806.49,-1843.9,-987.90,-14925.,-93.168,-18549.,-6004.0,-3869.3,-2155.2,66.383,2364.8,2156.3,895.93,320.22,1652.0,1686.6,0.0000,5801.9,4449.7,4252.8,3658.0,0.0000,-352.41,-106.73,-63.286,-44.256,-33.267,-587.69,0.0000,-1039.9,-1507.5,-739.88,-1165.5
1686.000000000,86.589,1988.9,2027.1,838.01,285.81,1531.5,967.16,3.8954,4745.5,2746.8,3370.4,2088.9,0.0000,-5990.5,-6606.7,-805.52,-1843.9,-984.94,-14923.,-93.141,-18547.,-6003.6,-3868.9,-2154.8,66.184,2357.8,2149.9,893.19,319.13,1647.1,1686.6,0.0000,5799.0,4449.7,4252.8,3658.0,0.0000,-351.39,-106.44,-63.090,-44.123,-33.130,-587.69,0.0000,-1039.8,-1507.5,-739.85,-1165.4
1687.000000000,86.784,1989.8,2030.8,837.13,285.71,1528.4,967.16,3.8957,4743.5,2746.8,3370.4,2088.9,0.0000,-5994.5,-6609.1,-804.48,-1843.9,-982.00,-14922.,-93.112,-18545.,-6003.3,-3868.5,-2154.3,65.930,2348.7,2141.6,890.15,317.87,1642.1,1686.6,0.0000,5796.0,4449.7,4252.8,3658.0,0.0000,-350.08,-106.07,-62.855,-43.953,-32.990,-587.69,0.0000,-1039.8,-1507.4,-739.82,-1165.3
1688.000000000,86.634,1988.1,2028.5,836.86,284.90,1525.1,967.16,3.8960,4741.4,2746.8,3370.4,2089.0,0.0000,-5997.7,-6611.1,-803.38,-1843.7,-979.03,-14920.,-93.084,-18543.,-6002.9,-3868.1,-2153.9,65.654,2338.9,2132.7,887.06,316.55,1637.2,1686.6,0.0000,5793.0,4449.7,4252.8,3658.0,0.0000,-348.64,-105.65,-62.608,-43.769,-32.853,-587.69,0.0000,-1039.8,-1507.4,-739.79,-1165.2
1689.000000000,86.419,1984.5,2027.7,836.67,283.96,1521.7,967.16,3.8962,4739.2,2746.9,3370.3,2089.0,0.0000,-6000.4,-6612.7,-802.22,-1843.4,-976.05,-14918.,-93.056,-18541.,-6002.6,-3867.7,-2153.4,65.456,2331.8,2126.2,884.91,315.60,1633.8,1686.6,0.0000,5791.1,4449.7,4252.8,3658.0,0.0000,-347.61,-105.36,-62.430,-43.637,-32.750,-587.69,0.0000,-1039.8,-1507.3,-739.76,-1165.2
1690.000000000,86.199,1981.4,2028.1,834.84,283.08,1518.2,967.16,3.7513,4736.9,2746.9,3370.3,2089.1,0.0000,-6002.7,-6613.9,-801.04,-1843.1,-973.07,-14916.,-93.027,-18540.,-6002.3,-3867.3,-2152.9,65.280,2325.6,2120.5,882.32,314.75,1629.1,1686.6,0.0000,5788.2,4449.7,4252.8,3658.0,0.0000,-346.70,-105.09,-62.251,-43.520,-32.616,-587.69,0.0000,-1039.8,-1507.2,-739.74,-1165.1
1691.000000000,85.820,1980.2,2026.9,833.53,282.12,1514.9,967.16,3.2816,4734.9,2747.0,3370.5,2089.1,0.0000,-6004.6,-6614.9,-799.86,-1842.7,-970.07,-14915.,-92.999,-18538.,-6001.9,-3866.9,-2152.5,64.971,2314.6,2110.5,879.07,313.28,1624.1,1686.6,0.0000,5785.2,4449.7,4252.8,3658.0,0.0000,-345.08,-104.61,-61.981,-43.314,-32.488,-587.69,0.0000,-1039.7,-1507.2,-739.71,-1165.0
1692.000000000,85.454,1973.8,2020.9,833.91,281.00,1511.0,967.16,3.2819,4732.7,2747.0,3370.5,2089.2,0.0000,-6005.9,-6615.5,-798.66,-1842.3,-967.08,-14913.,-92.971,-18536.,-6001.6,-3866.5,-2152.0,64.663,2303.6,2100.5,875.85,311.81,1619.2,1686.6,0.0000,5782.3,4449.7,4252.8,3658.0,0.0000,-343.45,-104.12,-61.713,-43.109,-32.366,-587.69,0.0000,-1039.7,-1507.1,-739.68,-1164.9
1693.000000000,85.184,1968.0,2012.8,833.05,279.88,1507.1,967.17,3.2822,4730.4,2746.8,3370.5,2089.3,0.0000,-6006.6,-6615.8,-797.45,-1841.9,-964.09,-14911.,-92.942,-18534.,-6001.2,-3866.1,-2151.6,64.347,2292.3,2090.2,872.55,310.30,1614.2,1686.6,0.0000,5779.3,4449.7,4252.8,3658.0,0.0000,-341.77,-103.61,-61.437,-42.898,-32.242,-587.69,0.0000,-1039.7,-1507.1,-739.65,-1164.8
1694.000000000,84.895,1963.0,2006.6,830.75,278.67,1503.2,967.17,3.2825,4728.8,2746.8,3370.5,2089.4,0.0000,-6006.6,-6615.8,-796.21,-1841.4,-961.10,-14909.,-92.914,-18532.,-6000.9,-3865.7,-2151.1,64.035,2281.2,2080.1,869.28,308.81,1609.3,1686.6,0.0000,5776.4,4449.7,4252.8,3658.0,0.0000,-340.11,-103.11,-61.165,-42.690,-32.118,-587.69,0.0000,-1039.7,-1507.0,-739.62,-1164.7
1695.000000000,84.583,1954.9,2000.2,828.41,277.40,1499.6,967.17,3.2828,4727.5,2746.9,3370.5,2089.5,0.0000,-6006.2,-6615.7,-794.95,-1840.9,-958.09,-14907.,-92.885,-18530.,-6000.5,-3865.3,-2150.7,63.733,2270.4,2070.3,866.12,307.37,1604.5,1686.6,0.0000,5773.5,4449.7,4252.8,3658.0,0.0000,-338.50,-102.62,-60.901,-42.489,-31.998,-587.69,0.0000,-1039.7,-1507.0,-739.59,-1164.6
1696.000000000,84.275,1947.1,1993.2,825.76,276.14,1496.3,967.17,3.2830,4725.7,2746.9,3370.6,2089.6,0.0000,-6005.4,-6615.4,-793.67,-1840.4,-955.08,-14906.,-92.856,-18528.,-6000.2,-3864.9,-2150.2,63.427,2259.5,2060.3,862.90,305.91,1599.5,1686.6,0.0000,5770.6,4449.7,4252.8,3658.0,0.0000,-336.85,-102.13,-60.634,-42.285,-31.876,-587.69,0.0000,-1039.6,-1506.9,-739.57,-1164.5
1697.000000000,83.967,1940.9,1988.5,823.00,275.07,1493.0,967.17,3.2833,4724.0,2747.0,3370.7,2089.6,0.0000,-6004.5,-6615.0,-792.38,-1839.9,-952.06,-14904.,-92.828,-18526.,-5999.8,-3864.5,-2149.7,136.16,2258.5,2078.7,862.77,306.29,1599.5,1686.6,0.0000,5770.6,4449.7,4252.8,3658.0,0.0000,-336.68,-102.49,-60.610,-42.268,-31.856,-587.69,0.0000,-1039.6,-1506.9,-739.54,-1164.4
1698.000000000,83.792,1936.5,1985.0,820.37,274.48,1490.0,967.17,3.2836,4721.9,2746.9,3370.7,2089.7,0.0000,-6003.7,-6614.5,-791.11,-1839.3,-949.06,-14902.,-92.801,-18524.,-5999.5,-3864.1,-2149.3,76.222,2255.2,2057.3,865.00,310.16,1604.7,1686.6,0.40729,5774.5,4450.3,4253.0,3658.5,0.0000,-336.15,-101.94,-60.592,-42.232,-31.927,-587.69,-0.18596E-01,-1039.6,-1506.8,-739.51,-1164.3
1699.000000000,83.640,1934.3,1980.6,818.37,273.77,1486.8,967.17,3.2839,4720.0,2746.7,3370.8,2089.7,0.0000,-6002.8,-6614.0,-789.84,-1838.8,-946.07,-14900.,-92.774,-18522.,-5999.1,-3863.7,-2148.8,63.127,2248.9,2050.6,862.21,304.52,1601.1,1686.6,0.0000,5771.6,4449.7,4252.8,3658.0,0.0000,-335.19,-101.62,-60.440,-42.085,-31.851,-587.69,0.0000,-1039.6,-1506.8,-739.48,-1164.2
1700.000000000,83.470,1930.5,1975.9,816.79,273.33,1483.9,967.17,3.2842,4717.9,2746.5,3370.9,2089.8,0.0000,-6001.7,-6613.4,-788.58,-1838.2,-943.11,-14899.,-92.746,-18520.,-5998.8,-3863.3,-2148.4,74.601,2314.1,2118.6,864.39,304.72,1602.9,1686.6,0.0000,5774.1,4449.7,4252.9,3658.0,0.0000,-335.48,-103.10,-60.476,-42.112,-31.857,-587.69,0.0000,-1039.6,-1506.7,-739.45,-1164.2
1701.000000000,83.436,1927.6,1972.4,815.38,273.13,1481.3,967.17,3.2845,4716.0,2746.5,3370.9,2090.0,0.0000,-6000.6,-6612.8,-787.32,-1837.7,-940.17,-14897.,-92.719,-18518.,-5998.4,-3862.9,-2147.9,62.950,2242.6,2044.9,860.40,303.68,1598.4,1686.6,0.0000,5770.0,4449.7,4252.8,3658.0,0.0000,-334.20,-101.32,-60.281,-41.967,-31.755,-587.69,0.0000,-1039.5,-1506.6,-739.42,-1164.1
1702.000000000,83.298,1922.6,1967.8,814.69,272.37,1478.7,967.17,3.2848,4714.4,2746.6,3371.0,2090.1,0.0000,-5999.2,-6612.1,-786.06,-1837.1,-937.27,-14895.,-92.691,-18516.,-5998.1,-3862.5,-2147.5,62.713,2234.1,2037.2,857.76,302.55,1594.3,1686.6,0.0000,5767.5,4449.7,4252.8,3658.0,0.0000,-332.90,-100.93,-60.068,-41.809,-31.649,-587.69,0.0000,-1039.5,-1506.6,-739.40,-1164.0
1703.000000000,83.131,1916.5,1961.7,813.77,271.61,1476.1,967.17,3.2851,4712.3,2746.6,3371.1,2090.2,0.0000,-5997.7,-6611.2,-784.79,-1836.6,-934.38,-14893.,-92.663,-18514.,-5997.7,-3862.1,-2147.0,62.478,2225.7,2029.5,855.18,301.42,1590.2,1686.6,0.0000,5765.1,4449.7,4252.8,3658.0,0.0000,-331.62,-100.54,-59.858,-41.652,-31.545,-587.69,0.0000,-1039.5,-1506.5,-739.37,-1163.9
1704.000000000,83.018,1910.7,1955.1,812.66,270.71,1473.3,967.17,3.2854,4710.3,2746.7,3371.0,2090.2,0.0000,-5995.8,-6610.1,-783.52,-1835.9,-931.49,-14891.,-92.635,-18512.,-5997.3,-3861.7,-2146.6,62.239,2217.2,2021.7,852.55,300.28,1586.1,1686.6,0.0000,5762.6,4449.7,4252.8,3658.0,0.0000,-330.31,-100.13,-59.644,-41.493,-31.440,-587.69,0.0000,-1039.5,-1506.5,-739.34,-1163.8
1705.000000000,82.783,1903.8,1949.0,811.74,269.72,1470.1,967.17,2.7890,4708.3,2747.0,3371.0,2090.3,0.0000,-5993.8,-6608.9,-782.24,-1835.3,-928.59,-14890.,-92.606,-18510.,-5997.0,-3861.4,-2146.1,61.967,2207.6,2012.9,849.52,298.98,1581.3,1686.6,0.0000,5759.8,4449.7,4252.8,3658.0,0.0000,-328.82,-99.680,-59.402,-41.312,-31.322,-587.69,0.0000,-1039.4,-1506.4,-739.31,-1163.7
1706.000000000,82.529,1896.8,1942.3,810.12,268.64,1466.8,967.17,2.6702,4706.4,2747.1,3371.0,2090.4,0.0000,-5991.5,-6607.5,-780.95,-1834.6,-925.68,-14888.,-92.578,-18508.,-5996.6,-3861.0,-2145.7,61.686,2197.5,2003.8,846.37,297.64,1576.3,1686.6,0.0000,5756.8,4449.7,4252.8,3658.0,0.0000,-327.28,-99.208,-59.150,-41.124,-31.199,-587.69,0.0000,-1039.4,-1506.4,-739.28,-1163.6
1707.000000000,82.240,1889.5,1938.4,808.19,267.51,1463.3,967.17,2.6705,4704.5,2747.2,3371.1,2090.5,0.0000,-5989.1,-6605.9,-779.66,-1833.9,-922.76,-14886.,-92.550,-18506.,-5996.3,-3860.6,-2145.2,61.400,2187.4,1994.5,843.16,296.27,1571.1,1686.6,0.0000,5753.8,4449.7,4252.8,3658.0,0.0000,-325.71,-98.727,-58.894,-40.934,-31.074,-587.69,0.0000,-1039.4,-1506.3,-739.25,-1163.5
1708.000000000,81.799,1882.2,1930.4,806.02,266.33,1459.9,967.17,2.6708,4702.4,2747.2,3371.1,2090.6,0.0000,-5986.5,-6604.2,-778.36,-1833.2,-919.83,-14884.,-92.521,-18504.,-5995.9,-3860.2,-2144.8,61.124,2177.5,1985.5,840.12,294.95,1566.3,1686.6,0.0000,5750.9,4449.7,4252.8,3658.0,0.0000,-324.19,-98.260,-58.648,-40.750,-30.955,-587.69,0.0000,-1039.4,-1506.3,-739.23,-1163.4
1709.000000000,81.536,1874.2,1922.4,803.76,265.18,1456.1,967.18,2.6712,4700.5,2747.3,3371.1,2090.7,0.0000,-5983.7,-6602.4,-777.05,-1832.5,-916.89,-14883.,-92.493,-18502.,-5995.5,-3859.8,-2144.3,60.846,2167.6,1976.5,836.97,293.62,1561.3,1686.6,0.0000,5747.9,4449.7,4252.8,3658.0,0.0000,-322.65,-97.788,-58.398,-40.564,-30.832,-587.69,0.0000,-1039.4,-1506.2,-739.20,-1163.3
1710.000000000,81.256,1866.0,1915.4,802.43,264.02,1452.4,967.18,2.6715,4698.9,2747.0,3371.2,2090.8,0.0000,-5980.7,-6600.5,-775.73,-1831.7,-913.96,-14881.,-92.465,-18501.,-5995.2,-3859.4,-2143.9,60.569,2157.7,1967.5,833.81,292.29,1556.2,1686.6,0.0000,5744.9,4449.7,4252.8,3658.0,0.0000,-321.12,-97.316,-58.148,-40.379,-30.708,-587.69,0.0000,-1039.3,-1506.2,-739.17,-1163.2
1711.000000000,80.976,1858.2,1909.5,800.08,262.90,1448.8,967.17,2.6718,4697.2,2747.1,3371.2,2090.9,0.0000,-5977.6,-6598.5,-774.39,-1831.0,-911.03,-14879.,-92.436,-18499.,-5994.8,-3859.0,-2143.4,60.315,2148.7,1959.3,830.91,291.08,1551.5,1686.6,0.0000,5742.1,4449.7,4252.8,3658.0,0.0000,-319.71,-96.880,-57.918,-40.210,-30.592,-587.69,0.0000,-1039.3,-1506.1,-739.14,-1163.1
1712.000000000,80.709,1850.6,1902.3,797.40,261.84,1445.4,967.13,2.6722,4695.6,2747.1,3371.2,2091.0,0.0000,-5974.3,-6596.4,-773.04,-1830.2,-908.08,-14877.,-92.408,-18497.,-5994.5,-3858.6,-2143.0,60.068,2139.9,1951.2,828.08,289.90,1547.0,1686.6,0.0000,5739.3,4449.7,4252.8,3658.0,0.0000,-318.33,-96.455,-57.694,-40.045,-30.479,-587.69,0.0000,-1039.3,-1506.0,-739.11,-1163.1
1713.000000000,80.450,1843.0,1894.8,794.78,260.79,1442.0,967.10,2.6725,4694.0,2747.2,3371.2,2091.0,0.0000,-5970.9,-6594.3,-771.69,-1829.4,-905.13,-14876.,-92.380,-18495.,-5994.1,-3858.2,-2142.5,59.826,2131.3,1943.4,825.29,288.74,1542.5,1686.6,0.0000,5736.6,4449.7,4252.8,3658.0,0.0000,-316.97,-96.037,-57.474,-39.884,-30.367,-587.69,0.0000,-1039.3,-1506.0,-739.08,-1163.0
1714.000000000,80.196,1835.9,1887.8,792.15,259.76,1439.2,967.10,2.6728,4692.3,2747.1,3371.2,2091.0,0.0000,-5967.3,-6592.1,-770.33,-1828.6,-902.16,-14874.,-92.351,-18493.,-5993.8,-3857.8,-2142.1,59.579,2122.5,1935.4,822.43,287.56,1537.8,1686.6,0.0000,5733.9,4449.7,4252.8,3658.0,0.0000,-315.59,-95.611,-57.250,-39.720,-30.252,-587.69,0.0000,-1039.3,-1505.9,-739.06,-1162.9
1715.000000000,79.997,1828.9,1880.4,789.50,258.76,1435.6,967.10,2.6731,4690.3,2747.0,3371.2,2091.2,0.0000,-5963.5,-6589.9,-768.96,-1827.7,-899.21,-14872.,-92.323,-18491.,-5993.4,-3857.4,-2141.7,59.339,2113.9,1927.5,819.63,286.41,1533.3,1686.6,0.0000,5731.1,4449.7,4252.8,3658.0,0.0000,-314.24,-95.195,-57.030,-39.559,-30.138,-587.69,0.0000,-1039.2,-1505.9,-739.03,-1162.8
1716.000000000,79.897,1821.8,1873.2,786.90,257.79,1431.9,967.10,2.6734,4688.3,2747.0,3371.2,2091.3,0.0000,-5959.6,-6587.6,-767.59,-1826.9,-896.24,-14870.,-92.295,-18489.,-5993.1,-3857.0,-2141.2,59.102,2105.5,1919.8,816.84,285.27,1528.7,1686.6,0.0000,5728.4,4449.7,4252.8,3658.0,0.0000,-312.90,-94.784,-56.814,-39.401,-30.026,-587.69,0.0000,-1039.2,-1505.8,-739.00,-1162.7
1717.000000000,79.661,1814.7,1866.1,784.24,256.81,1428.0,967.10,2.6721,4686.1,2747.1,3371.2,2091.5,0.0000,-5955.5,-6585.3,-766.21,-1826.1,-893.28,-14869.,-92.267,-18487.,-5992.7,-3856.6,-2140.8,58.861,2096.9,1912.0,814.00,284.12,1524.0,1686.6,0.0000,5725.6,4449.7,4252.8,3658.0,0.0000,-311.55,-94.365,-56.593,-39.241,-29.910,-587.69,0.0000,-1039.2,-1505.8,-738.97,-1162.6
1718.000000000,79.439,1807.4,1858.6,781.73,255.80,1423.9,967.10,2.6663,4683.7,2747.1,3371.3,2091.5,0.0000,-5951.4,-6582.9,-764.83,-1825.2,-890.32,-14867.,-92.239,-18485.,-5992.4,-3856.2,-2140.3,58.606,2087.8,1903.7,810.95,282.89,1519.0,1686.6,0.0000,5722.6,4449.7,4252.8,3658.0,0.0000,-310.11,-93.923,-56.358,-39.070,-29.788,-587.69,0.0000,-1039.2,-1505.7,-738.94,-1162.5
1719.000000000,79.290,1800.0,1850.8,779.18,254.77,1419.7,967.10,2.6666,4681.1,2747.2,3371.3,2091.6,0.0000,-5947.0,-6580.5,-763.44,-1824.4,-887.35,-14865.,-92.210,-18483.,-5992.0,-3855.8,-2139.9,58.341,2078.4,1895.1,807.78,281.62,1513.7,1686.6,0.0000,5719.5,4449.7,4252.8,3658.0,0.0000,-308.62,-93.466,-56.114,-38.894,-29.661,-587.69,0.0000,-1039.2,-1505.7,-738.92,-1162.4
1720.000000000,79.082,1792.4,1842.8,776.62,253.73,1415.7,967.10,2.6669,4678.6,2747.2,3371.4,2091.7,0.0000,-5942.5,-6578.0,-762.05,-1823.5,-884.38,-14863.,-92.182,-18481.,-5991.7,-3855.5,-2139.4,58.087,2069.3,1886.9,804.72,280.40,1508.7,1686.6,0.0000,5716.4,4449.7,4252.8,3658.0,0.0000,-307.19,-93.024,-55.879,-38.725,-29.538,-587.69,0.0000,-1039.1,-1505.6,-738.89,-1162.3
1721.000000000,78.974,1784.8,1835.0,773.97,252.69,1411.8,967.06,2.6672,4676.0,2747.3,3371.4,2091.7,0.0000,-5937.9,-6575.4,-760.65,-1822.6,-881.41,-14862.,-92.154,-18479.,-5991.3,-3855.1,-2139.0,57.837,2060.4,1878.8,801.68,279.20,1503.6,1686.6,0.0000,5713.4,4449.7,4252.8,3658.0,0.0000,-305.77,-92.589,-55.648,-38.558,-29.415,-587.69,0.0000,-1039.1,-1505.6,-738.86,-1162.2
1722.000000000,78.687,1777.2,1827.2,771.34,251.64,1407.5,967.06,2.6675,4673.6,2747.4,3371.5,2091.8,0.0000,-5933.2,-6572.8,-759.24,-1821.7,-878.43,-14860.,-92.126,-18478.,-5991.0,-3854.7,-2138.6,57.599,2052.0,1871.0,798.78,278.06,1498.7,1686.6,0.0000,5710.5,4449.7,4252.8,3658.0,0.0000,-304.43,-92.173,-55.427,-38.400,-29.296,-587.69,0.0000,-1039.1,-1505.5,-738.83,-1162.2
1723.000000000,78.281,1770.0,1819.9,768.68,250.64,1403.0,967.03,2.6678,4671.4,2747.4,3371.7,2091.9,0.0000,-5928.4,-6570.2,-757.84,-1820.8,-875.45,-14858.,-92.098,-18476.,-5990.6,-3854.3,-2138.1,57.361,2043.4,1863.3,795.85,276.92,1493.8,1686.6,0.0000,5707.5,4449.7,4252.8,3658.0,0.0000,-303.07,-91.755,-55.204,-38.241,-29.176,-587.69,0.0000,-1039.1,-1505.5,-738.80,-1162.1
1724.000000000,78.037,1763.0,1812.6,766.08,249.65,1398.7,967.03,2.6682,4669.0,2747.5,3371.8,2091.9,0.0000,-5923.5,-6567.6,-756.43,-1819.9,-872.46,-14856.,-92.070,-18474.,-5990.3,-3853.9,-2137.7,57.141,2035.6,1856.2,793.23,275.87,1489.5,1686.6,0.0000,5705.0,4449.7,4252.8,3658.0,0.0000,-301.82,-91.368,-55.002,-38.094,-29.069,-587.69,0.0000,-1039.0,-1505.4,-738.77,-1162.0
1725.000000000,77.802,1756.2,1805.5,763.46,248.69,1394.5,967.03,2.6685,4666.5,2747.5,3371.8,2092.0,0.0000,-5918.5,-6565.0,-755.02,-1818.9,-869.47,-14855.,-92.042,-18472.,-5989.9,-3853.5,-2137.3,56.904,2027.2,1848.5,790.29,274.73,1484.5,1686.6,0.0000,5702.0,4449.7,4252.8,3658.0,0.0000,-300.47,-90.952,-54.780,-37.936,-28.948,-587.69,0.0000,-1039.0,-1505.4,-738.75,-1161.9
1726.000000000,77.569,1749.2,1798.6,760.87,247.72,1390.3,967.03,2.6688,4664.1,2747.6,3372.0,2092.1,0.0000,-5913.5,-6562.4,-753.61,-1818.0,-866.48,-14853.,-92.014,-18470.,-5989.6,-3853.1,-2136.8,56.673,2018.9,1840.9,787.39,273.61,1479.6,1686.6,0.0000,5699.0,4449.7,4252.8,3658.0,0.0000,-299.14,-90.545,-54.563,-37.782,-28.829,-587.69,0.0000,-1039.0,-1505.3,-738.72,-1161.8
1727.000000000,77.234,1742.2,1791.5,758.26,246.78,1386.2,967.03,2.6691,4661.6,2747.6,3372.1,2092.1,0.0000,-5908.3,-6559.7,-752.19,-1817.1,-863.50,-14851.,-91.986,-18468.,-5989.2,-3852.8,-2136.4,56.451,2011.0,1833.7,784.83,272.55,1475.4,1686.6,0.0000,5696.6,4449.7,4252.8,3658.0,0.0000,-297.88,-90.154,-54.361,-37.634,-28.725,-587.69,0.0000,-1039.0,-1505.3,-738.69,-1161.7
1728.000000000,76.950,1735.4,1784.6,755.68,245.86,1381.9,967.03,2.6694,4659.1,2747.7,3372.2,2092.2,0.0000,-5903.1,-6557.0,-750.78,-1816.1,-860.52,-14849.,-91.958,-18466.,-5988.9,-3852.4,-2136.0,56.235,2003.3,1826.7,782.08,271.51,1470.7,1686.6,0.0000,5693.7,4449.7,4252.8,3658.0,0.0000,-296.63,-89.771,-54.156,-37.490,-28.610,-587.69,0.0000,-1039.0,-1505.2,-738.66,-1161.6
1729.000000000,76.699,1733.4,1781.7,753.09,245.65,1377.9,967.03,2.6697,4656.6,2747.7,3372.3,2092.3,0.0000,-5898.2,-6554.5,-749.41,-1815.2,-857.55,-14848.,-91.932,-18464.,-5988.5,-3852.0,-2135.6,79.372,2043.8,1877.6,794.74,277.23,1491.7,1686.6,1.1597,5707.0,4450.7,4253.2,3658.5,0.0000,-301.39,-91.654,-55.004,-38.110,-29.007,-587.69,-0.52952E-01,-1039.0,-1505.1,-738.64,-1161.5
1730.000000000,76.849,1745.0,1789.4,750.96,247.54,1374.9,967.02,2.6714,4654.3,2747.8,3372.4,2092.4,0.0000,-5894.3,-6552.7,-748.12,-1814.5,-854.60,-14846.,-91.907,-18462.,-5988.2,-3851.6,-2135.2,143.93,2165.5,2022.2,816.74,293.32,1519.1,1686.6,69.372,5728.5,4463.0,4266.3,3671.5,0.0000,-305.95,-95.485,-55.743,-38.754,-29.344,-587.69,-3.1674,-1039.1,-1505.1,-738.67,-1161.6
1731.000000000,77.313,1776.8,1817.8,750.88,251.92,1374.7,967.02,2.7211,4652.7,2747.8,3372.4,2092.4,0.0000,-5892.6,-6552.4,-747.11,-1813.9,-851.78,-14844.,-91.885,-18460.,-5987.9,-3851.2,-2134.8,717.82,3374.6,3017.5,916.63,340.28,1687.3,1687.0,1030.0,5840.6,4489.6,4293.1,3698.3,0.0000,-330.24,-120.61,-60.306,-41.790,-32.343,-587.69,-47.027,-1039.5,-1505.0,-738.77,-1161.9
1732.000000000,79.343,1861.7,1892.3,775.60,265.71,1461.4,966.99,2.7271,4663.7,2747.9,3372.4,2092.5,0.0000,-5896.1,-6555.5,-749.10,-1814.1,-852.10,-14842.,-91.866,-18458.,-5987.5,-3850.8,-2134.4,2021.8,4355.6,3962.7,2396.7,485.39,5059.7,1701.8,1444.6,7992.7,4644.0,4426.9,3827.5,0.0000,-365.35,-146.65,-103.17,-46.663,-99.323,-587.90,-65.961,-1042.4,-1505.0,-739.39,-1163.5
1733.000000000,83.840,1978.6,1997.3,935.46,281.47,1804.2,966.98,2.7275,4759.2,2747.9,3372.6,2092.6,0.0000,-5906.0,-6562.8,-755.18,-1815.0,-859.87,-14841.,-91.848,-18457.,-5987.2,-3850.4,-2134.0,385.41,3132.6,2740.2,2416.2,561.79,5100.9,1758.3,993.14,8011.0,4696.5,4486.0,3887.7,0.0000,-374.52,-122.56,-104.61,-48.468,-99.642,-588.69,-45.346,-1042.6,-1504.9,-739.64,-1164.3
1734.000000000,86.739,2059.3,2081.2,1211.4,309.53,2270.0,966.98,2.7278,4866.0,2748.0,3373.2,2092.9,0.0000,-5918.9,-6571.9,-760.59,-1816.1,-875.60,-14839.,-91.827,-18459.,-5986.9,-3850.1,-2133.6,183.80,2773.4,2522.8,2336.8,476.59,5014.4,1855.1,209.16,7990.7,4599.3,4485.5,3888.8,0.0000,-382.35,-119.46,-105.72,-48.950,-99.421,-590.05,-9.5501,-1042.3,-1504.9,-739.61,-1164.2
1735.000000000,89.966,2112.3,2136.4,1423.8,326.10,2635.6,966.99,2.7282,5015.0,2748.0,3374.4,2093.7,0.0000,-5932.9,-6580.9,-768.27,-1817.2,-900.02,-14837.,-91.805,-18459.,-5986.5,-3849.7,-2133.2,72.861,2595.6,2366.8,2248.3,401.40,4904.8,1712.4,0.0000,7779.9,4486.1,4285.3,3690.1,0.0000,-384.48,-116.64,-106.11,-48.760,-99.219,-588.05,0.0000,-1039.4,-1504.9,-738.62,-1161.5
1736.000000000,92.001,2139.4,2169.6,1613.9,330.87,2866.4,966.99,16.859,5107.8,2747.9,3374.4,2093.3,0.0000,-5946.6,-6589.2,-776.74,-1818.1,-918.83,-14836.,-91.781,-18460.,-5986.2,-3849.3,-2132.8,72.774,2592.5,2364.0,2184.0,393.55,4873.9,1708.2,0.0000,7773.2,4473.6,4278.1,3682.2,0.0000,-384.19,-116.62,-106.15,-48.656,-99.395,-587.99,0.0000,-1039.3,-1504.8,-738.56,-1161.3
1737.000000000,92.628,2151.4,2184.0,1754.8,332.48,3032.1,966.99,26.394,5175.3,2748.6,3375.4,2093.4,0.0000,-5959.0,-6596.5,-785.91,-1818.8,-933.99,-14834.,-91.756,-18461.,-5985.9,-3848.9,-2132.4,72.549,2584.5,2356.7,2165.9,379.37,4857.0,1705.6,0.0000,7754.5,4457.4,4261.1,3665.8,0.0000,-383.19,-116.37,-106.10,-48.425,-99.617,-587.95,0.0000,-1039.0,-1504.8,-738.45,-1161.0
1738.000000000,93.732,2159.6,2194.2,1837.8,332.73,3165.1,966.99,35.876,5308.5,2749.7,3377.1,2093.9,0.0000,-5970.5,-6603.0,-798.96,-1819.3,-947.06,-14833.,-91.732,-18461.,-5985.5,-3848.6,-2132.0,72.664,2897.3,2463.9,2368.3,486.69,5052.7,1713.2,600.93,7954.4,4650.3,4453.5,3857.7,0.0000,-384.44,-118.87,-106.30,-49.160,-100.76,-588.06,-27.438,-1041.7,-1504.7,-739.35,-1163.4
1739.000000000,93.872,2164.2,2205.9,1914.3,332.66,3219.1,966.99,26.741,5419.5,2750.2,3376.4,2093.8,0.0000,-5981.2,-6608.7,-809.54,-1819.7,-958.67,-14831.,-91.707,-18462.,-5985.2,-3848.2,-2131.6,72.502,2582.9,2355.1,2157.0,371.43,4848.8,1701.3,0.0000,7751.6,4455.4,4258.0,3662.0,0.0000,-383.28,-116.50,-106.30,-48.346,-100.13,-587.89,0.0000,-1038.9,-1504.7,-738.38,-1160.8
1740.000000000,93.530,2172.1,2216.4,1924.5,331.92,3391.2,966.99,28.756,5701.5,2750.1,3376.2,2094.1,0.0000,-5991.1,-6614.1,-818.33,-1820.0,-969.25,-14830.,-91.682,-18464.,-5984.9,-3847.8,-2131.2,72.208,2572.4,2345.6,2152.8,368.76,4846.2,1699.7,0.0000,7745.9,4454.7,4256.3,3661.5,0.0000,-381.89,-116.11,-106.20,-48.142,-100.36,-587.87,0.0000,-1038.8,-1504.6,-738.35,-1160.7
1741.000000000,93.187,2171.6,2214.6,1931.4,331.16,3668.3,966.99,31.591,5947.9,2751.6,3375.8,2094.2,0.0000,-5999.8,-6618.7,-826.08,-1820.2,-979.11,-14829.,-91.657,-18466.,-5984.6,-3847.5,-2130.8,71.882,2560.8,2335.0,2148.1,366.73,4842.9,1698.4,0.0000,7741.5,4450.3,4253.1,3658.3,0.0000,-380.32,-115.66,-106.07,-47.921,-100.58,-587.85,0.0000,-1038.7,-1504.6,-738.31,-1160.5
1742.000000000,92.824,2167.2,2208.6,1934.0,330.05,3949.9,967.00,36.778,6109.9,2755.0,3378.0,2094.9,0.0000,-6007.2,-6622.6,-833.15,-1820.4,-988.45,-14827.,-91.631,-18468.,-5984.4,-3847.1,-2130.4,71.559,2549.3,2324.5,2146.3,365.22,4842.4,1697.3,0.0000,7740.9,4449.7,4252.8,3658.0,0.0000,-378.75,-115.21,-105.94,-47.706,-100.80,-587.84,0.0000,-1038.7,-1504.5,-738.28,-1160.4
1743.000000000,92.473,2167.1,2202.0,1945.8,328.79,4045.0,967.00,34.072,6212.7,2756.9,3376.7,2095.7,0.0000,-6013.4,-6626.0,-839.74,-1820.5,-997.42,-14826.,-91.605,-18471.,-5984.2,-3846.8,-2130.0,71.220,2537.2,2313.5,2144.8,363.64,4842.3,1696.6,0.0000,7740.9,4449.7,4252.8,3658.0,0.0000,-377.08,-114.72,-105.79,-47.480,-101.01,-587.83,0.0000,-1038.7,-1504.5,-738.26,-1160.4
1744.000000000,92.044,2161.8,2199.4,1984.4,327.55,4085.4,967.00,35.377,6250.2,2756.2,3376.1,2096.6,0.0000,-6018.5,-6629.1,-845.93,-1820.6,-1006.1,-14825.,-91.580,-18474.,-5984.0,-3846.4,-2129.5,70.988,2542.1,2305.9,2243.3,362.55,4842.2,1695.7,691.88,7953.4,4652.4,4252.8,3664.8,0.0000,-375.98,-114.40,-105.70,-47.325,-101.22,-587.82,-31.590,-1041.6,-1504.4,-738.24,-1160.4
1745.000000000,91.879,2157.0,2195.0,1999.0,326.68,4088.1,967.01,31.600,6271.4,2753.6,3375.5,2097.5,0.0000,-6022.9,-6632.0,-851.80,-1820.7,-1014.7,-14825.,-91.555,-18477.,-5983.8,-3846.1,-2129.1,70.728,2519.7,2297.5,2142.6,361.34,4842.2,1695.0,0.0000,7740.9,4449.7,4252.8,3658.0,0.0000,-374.69,-114.03,-105.60,-47.152,-101.50,-587.81,0.0000,-1038.6,-1504.4,-738.22,-1160.2
1746.000000000,91.597,2152.9,2191.1,1997.8,325.60,4098.7,966.98,36.492,6270.8,2753.1,3374.6,2097.1,0.0000,-6027.1,-6634.5,-857.37,-1820.7,-1023.1,-14824.,-91.529,-18480.,-5983.6,-3845.8,-2128.7,70.405,2508.2,2287.0,2141.2,359.83,4842.0,1694.4,0.0000,7740.9,4449.7,4252.8,3658.0,0.0000,-373.07,-113.55,-105.45,-46.937,-101.81,-587.80,0.0000,-1038.6,-1504.3,-738.19,-1160.1
1747.000000000,91.240,2145.2,2188.9,1996.7,324.43,4126.8,966.97,37.840,6273.1,2752.6,3374.0,2096.4,0.0000,-6031.2,-6636.7,-862.66,-1820.6,-1031.9,-14823.,-91.504,-18482.,-5983.4,-3845.5,-2128.3,70.073,2496.3,2276.2,2139.7,358.28,4841.9,1693.8,0.0000,7740.9,4449.7,4252.8,3658.0,0.0000,-371.39,-113.05,-105.28,-46.715,-102.10,-587.79,0.0000,-1038.6,-1504.3,-738.17,-1160.0
1748.000000000,90.899,2139.0,2180.5,1995.5,323.13,4161.1,966.97,35.926,6306.3,2752.4,3373.7,2096.9,0.0000,-6034.6,-6638.5,-867.71,-1820.6,-1041.1,-14822.,-91.478,-18485.,-5983.2,-3845.1,-2128.0,69.727,2484.0,2265.0,2138.1,356.67,4841.8,1693.4,0.0000,7740.9,4449.7,4252.8,3658.0,0.0000,-369.63,-112.52,-105.11,-46.485,-102.40,-587.78,0.0000,-1038.6,-1504.2,-738.15,-1159.9
1749.000000000,90.728,2131.0,2171.0,1994.2,321.68,4224.9,966.99,35.193,6336.1,2751.5,3373.6,2097.1,0.0000,-6037.3,-6640.0,-872.51,-1820.4,-1050.5,-14821.,-91.452,-18488.,-5982.9,-3844.8,-2127.6,69.394,2472.1,2254.2,2136.6,355.11,4841.7,1693.1,0.0000,7740.9,4449.7,4252.8,3658.0,0.0000,-367.93,-112.01,-104.94,-46.263,-102.68,-587.78,0.0000,-1038.6,-1504.2,-738.12,-1159.8
1750.000000000,90.401,2121.0,2161.6,2004.4,320.37,4241.5,966.99,31.092,6335.7,2752.1,3373.3,2097.1,0.0000,-6039.4,-6641.2,-877.10,-1820.2,-1059.8,-14821.,-91.426,-18491.,-5982.6,-3844.5,-2127.2,69.114,2462.1,2245.1,2135.4,353.80,4841.6,1692.7,0.0000,7740.9,4449.7,4252.8,3658.0,0.0000,-366.50,-111.58,-104.81,-46.076,-102.96,-587.77,0.0000,-1038.6,-1504.2,-738.10,-1159.7
1751.000000000,89.993,2112.3,2152.4,2014.1,319.17,4258.7,967.00,30.703,6335.6,2753.4,3373.3,2096.8,0.0000,-6041.1,-6642.1,-881.48,-1820.0,-1069.0,-14820.,-91.400,-18493.,-5982.4,-3844.1,-2126.8,68.836,2452.2,2236.0,2134.2,352.51,4841.5,1690.6,0.0000,7740.9,4449.7,4252.8,3658.0,0.0000,-365.08,-111.15,-104.67,-45.891,-103.23,-587.74,0.0000,-1038.6,-1504.1,-738.07,-1159.6
1752.000000000,89.694,2104.2,2144.2,2014.8,317.98,4257.8,967.00,31.440,6362.6,2755.3,3373.3,2096.8,0.0000,-6042.3,-6642.6,-885.67,-1819.7,-1077.9,-14819.,-91.374,-18496.,-5982.1,-3843.8,-2126.4,68.554,2442.2,2226.9,2132.9,351.19,4841.4,1687.7,0.0000,7740.9,4449.7,4252.8,3658.0,0.0000,-363.62,-110.70,-104.53,-45.702,-103.50,-587.70,0.0000,-1038.6,-1504.1,-738.05,-1159.5
1753.000000000,89.405,2098.2,2135.3,2014.1,316.82,4264.3,967.00,33.265,6378.8,2755.4,3373.4,2096.7,0.0000,-6043.1,-6642.9,-889.68,-1819.4,-1086.9,-14819.,-91.348,-18499.,-5981.8,-3843.5,-2126.0,68.264,2431.9,2217.5,2131.6,349.84,4841.3,1686.8,0.0000,7740.9,4449.7,4252.8,3658.0,0.0000,-362.11,-110.24,-104.38,-45.509,-103.76,-587.69,0.0000,-1038.6,-1504.0,-738.02,-1159.5
1754.000000000,89.223,2089.4,2127.3,2015.2,315.60,4281.5,967.00,36.140,6391.1,2756.3,3373.8,2097.3,0.0000,-6043.6,-6642.8,-893.53,-1819.1,-1096.2,-14818.,-91.322,-18501.,-5981.6,-3843.2,-2125.6,67.972,2421.5,2208.0,2130.3,348.48,4841.2,1686.6,0.0000,7740.9,4449.7,4252.8,3658.0,0.0000,-360.58,-109.77,-104.23,-45.315,-104.02,-587.69,0.0000,-1038.6,-1504.0,-738.00,-1159.4
1755.000000000,88.960,2080.6,2121.0,2014.1,314.39,4288.6,967.00,27.305,6400.2,2755.3,3373.6,2097.2,0.0000,-6043.7,-6642.5,-897.23,-1818.7,-1105.4,-14818.,-91.296,-18503.,-5981.4,-3842.9,-2125.2,67.672,2410.8,2198.2,2128.9,347.08,4841.1,1686.6,0.0000,7740.9,4449.7,4252.8,3658.0,0.0000,-359.00,-109.29,-104.07,-45.115,-104.27,-587.69,0.0000,-1038.6,-1503.9,-737.97,-1159.3
1756.000000000,88.407,2072.1,2121.5,2012.9,313.14,4294.2,967.01,25.672,6403.9,2753.3,3373.5,2097.2,0.0000,-6043.8,-6642.0,-900.78,-1818.3,-1114.3,-14817.,-91.270,-18506.,-5981.1,-3842.5,-2124.8,67.375,2400.2,2188.6,2127.6,345.69,4841.0,1686.6,0.0000,7740.9,4449.7,4252.8,3658.0,0.0000,-357.43,-108.80,-103.91,-44.916,-104.52,-587.69,0.0000,-1038.6,-1503.9,-737.95,-1159.2
1757.000000000,88.110,2065.1,2115.2,2011.7,311.96,4313.1,966.98,22.873,6420.9,2752.3,3373.3,2097.2,0.0000,-6043.8,-6641.2,-904.19,-1817.9,-1122.9,-14817.,-91.244,-18508.,-5980.8,-3842.2,-2124.4,67.103,2390.5,2179.8,2126.4,344.42,4840.9,1686.6,0.0000,7740.9,4449.7,4252.8,3658.0,0.0000,-355.99,-108.36,-103.77,-44.735,-104.76,-587.69,0.0000,-1038.6,-1503.8,-737.92,-1159.1
1758.000000000,87.800,2056.6,2106.6,2010.5,310.83,4330.4,966.97,27.516,6445.2,2753.3,3373.1,2097.3,0.0000,-6043.5,-6640.3,-907.47,-1817.5,-1131.0,-14817.,-91.217,-18510.,-5980.5,-3841.9,-2124.0,66.827,2380.7,2170.8,2125.2,343.13,4840.9,1686.6,0.0000,7740.9,4449.7,4252.8,3658.0,0.0000,-354.52,-107.90,-103.62,-44.551,-105.00,-587.69,0.0000,-1038.6,-1503.8,-737.89,-1159.0
1759.000000000,87.444,2048.2,2099.5,2011.3,309.72,4329.7,966.97,25.715,6476.7,2754.1,3373.2,2097.2,0.0000,-6043.1,-6639.3,-910.62,-1817.0,-1138.8,-14817.,-91.191,-18513.,-5980.2,-3841.6,-2123.6,66.579,2371.8,2162.7,2124.1,341.97,4840.8,1686.6,0.0000,7740.9,4449.7,4252.8,3658.0,0.0000,-353.19,-107.49,-103.49,-44.386,-105.23,-587.69,0.0000,-1038.6,-1503.7,-737.87,-1158.9
1760.000000000,87.179,2040.4,2097.0,2011.0,308.69,4341.9,966.97,18.943,6486.3,2755.1,3373.2,2097.3,0.0000,-6042.6,-6638.3,-913.67,-1816.5,-1146.4,-14816.,-91.165,-18515.,-5980.0,-3841.3,-2123.2,66.329,2362.9,2154.6,2122.9,340.81,4840.7,1686.6,0.0000,7740.9,4449.7,4252.8,3658.0,0.0000,-351.85,-107.07,-103.36,-44.220,-105.46,-587.69,0.0000,-1038.6,-1503.7,-737.84,-1158.8
1761.000000000,86.921,2032.7,2090.6,2009.9,307.66,4365.1,966.97,16.539,6502.4,2755.1,3373.2,2097.4,0.0000,-6041.9,-6637.0,-916.60,-1816.0,-1154.1,-14816.,-91.138,-18517.,-5979.7,-3841.0,-2122.8,66.066,2353.6,2146.1,2121.8,339.58,4840.6,1686.6,0.0000,7740.9,4449.7,4252.8,3658.0,0.0000,-350.44,-106.64,-103.22,-44.044,-105.68,-587.69,0.0000,-1038.6,-1503.6,-737.82,-1158.7
1762.000000000,86.533,2025.0,2082.6,2008.7,306.66,4382.2,966.97,18.911,6507.8,2754.9,3373.0,2097.6,0.0000,-6041.0,-6635.6,-919.43,-1815.5,-1163.4,-14816.,-91.112,-18519.,-5979.4,-3840.7,-2122.4,65.855,2346.1,2139.2,2120.8,338.60,4840.5,1686.6,0.0000,7740.9,4449.7,4252.8,3658.0,0.0000,-349.29,-106.28,-103.11,-43.904,-105.90,-587.69,0.0000,-1038.6,-1503.6,-737.79,-1158.6
1763.000000000,86.150,2017.6,2075.1,2007.7,305.76,4381.6,966.98,18.910,6507.6,2753.7,3373.2,2098.0,0.0000,-6039.9,-6634.1,-922.16,-1815.0,-1171.9,-14816.,-91.085,-18521.,-5979.1,-3840.5,-2122.0,65.645,2338.6,2132.4,2119.9,337.62,4840.5,1686.6,0.0000,7740.9,4449.7,4252.8,3658.0,0.0000,-348.15,-105.92,-103.00,-43.764,-106.11,-587.69,0.0000,-1038.6,-1503.5,-737.77,-1158.5
1764.000000000,85.924,2010.6,2067.9,2007.0,304.85,4382.3,966.98,14.045,6507.4,2752.7,3373.2,2098.1,0.0000,-6038.4,-6632.5,-924.80,-1814.5,-1179.6,-14816.,-91.059,-18522.,-5978.8,-3840.2,-2121.6,65.423,2330.7,2125.2,2118.9,336.58,4840.4,1686.6,0.0000,7740.9,4449.7,4252.8,3658.0,0.0000,-346.94,-105.55,-102.88,-43.615,-106.32,-587.69,0.0000,-1038.6,-1503.5,-737.74,-1158.4
1765.000000000,85.698,2003.9,2060.7,2005.8,303.95,4402.3,966.98,13.602,6507.2,2752.5,3373.2,2098.0,0.0000,-6036.8,-6630.9,-927.36,-1813.9,-1186.9,-14815.,-91.032,-18524.,-5978.5,-3839.9,-2121.2,65.184,2322.1,2117.4,2117.8,335.46,4840.3,1686.6,0.0000,7740.9,4449.7,4252.8,3658.0,0.0000,-345.63,-105.14,-102.75,-43.456,-106.53,-587.69,0.0000,-1038.7,-1503.4,-737.72,-1158.3
1766.000000000,85.422,1997.0,2053.3,2004.7,303.06,4409.2,966.98,13.602,6507.0,2752.9,3373.3,2097.9,0.0000,-6035.0,-6629.1,-929.83,-1813.3,-1193.9,-14815.,-91.006,-18526.,-5978.2,-3839.6,-2120.8,64.975,2314.7,2110.6,2116.9,334.49,4840.2,1686.6,0.0000,7740.9,4449.7,4252.8,3658.0,0.0000,-344.49,-104.78,-102.64,-43.317,-106.73,-587.69,0.0000,-1038.7,-1503.4,-737.69,-1158.2
1767.000000000,85.103,1990.2,2046.1,2003.7,302.19,4423.2,966.98,13.601,6506.8,2753.0,3373.4,2097.8,0.0000,-6033.0,-6627.3,-932.22,-1812.8,-1200.5,-14815.,-90.979,-18528.,-5977.9,-3839.3,-2120.4,64.733,2306.1,2102.8,2115.8,333.36,4840.2,1686.6,0.0000,7740.9,4449.7,4252.8,3658.0,0.0000,-343.16,-104.37,-102.51,-43.155,-106.94,-587.69,0.0000,-1038.7,-1503.3,-737.66,-1158.1
1768.000000000,84.870,1983.3,2038.1,2002.7,301.23,4427.6,966.98,13.601,6506.7,2754.0,3373.6,2097.9,0.0000,-6030.8,-6625.5,-934.53,-1812.2,-1206.9,-14815.,-90.952,-18530.,-5977.6,-3839.1,-2120.0,64.480,2297.1,2094.6,2114.7,332.18,4840.1,1686.6,0.0000,7740.9,4449.7,4252.8,3658.0,0.0000,-341.77,-103.94,-102.37,-42.987,-107.13,-587.69,0.0000,-1038.7,-1503.3,-737.64,-1158.0
1769.000000000,84.426,1975.7,2030.6,2001.6,300.27,4444.1,966.99,13.601,6506.5,2755.3,3373.8,2097.9,0.0000,-6028.3,-6623.6,-936.77,-1811.6,-1213.0,-14815.,-90.926,-18534.,-5977.3,-3838.8,-2119.6,64.234,2288.3,2086.6,2113.6,331.03,4840.0,1686.6,0.0000,7740.9,4449.7,4252.8,3658.0,0.0000,-340.41,-103.52,-102.23,-42.823,-107.33,-587.69,0.0000,-1038.7,-1503.2,-737.61,-1157.9
1770.000000000,84.158,1968.2,2022.9,2000.5,299.29,4443.6,966.99,13.599,6526.6,2754.6,3373.9,2097.9,0.0000,-6025.7,-6621.6,-938.93,-1810.9,-1219.0,-14814.,-90.899,-18537.,-5977.1,-3838.6,-2119.2,63.981,2279.3,2078.3,2112.4,329.85,4839.9,1686.6,0.0000,7740.9,4449.7,4252.8,3658.0,0.0000,-339.01,-103.09,-102.08,-42.654,-107.52,-587.69,0.0000,-1038.7,-1503.1,-737.59,-1157.9
1771.000000000,83.916,1960.9,2015.0,1999.5,298.30,4443.1,966.99,13.598,6528.2,2754.3,3374.1,2097.9,0.0000,-6022.9,-6619.5,-941.03,-1810.3,-1224.8,-14814.,-90.873,-18540.,-5976.8,-3838.3,-2118.8,63.736,2270.6,2070.4,2111.3,328.71,4839.8,1686.6,0.0000,7740.9,4449.7,4252.8,3658.0,0.0000,-337.66,-102.66,-101.94,-42.491,-107.70,-587.69,0.0000,-1038.7,-1503.1,-737.56,-1157.8
1772.000000000,83.667,1953.8,2006.9,1998.5,297.31,4444.8,966.99,13.598,6528.1,2753.5,3374.2,2098.1,0.0000,-6019.9,-6617.4,-943.07,-1809.6,-1230.4,-14814.,-90.846,-18542.,-5976.5,-3838.1,-2118.4,63.497,2262.0,2062.6,2110.3,327.59,4839.7,1686.6,0.0000,7740.9,4449.7,4252.8,3658.0,0.0000,-336.33,-102.25,-101.81,-42.331,-107.89,-587.69,0.0000,-1038.7,-1503.0,-737.54,-1157.7
1773.000000000,83.423,1946.7,1999.6,1997.4,296.35,4463.1,966.99,11.960,6538.0,2752.8,3374.2,2098.2,0.0000,-6016.7,-6615.2,-945.04,-1809.0,-1236.0,-14814.,-90.820,-18545.,-5976.2,-3837.8,-2118.0,63.281,2254.3,2055.6,2109.3,326.58,4839.7,1686.6,0.0000,7740.9,4449.7,4252.8,3658.0,0.0000,-335.12,-101.87,-101.69,-42.187,-108.07,-587.69,0.0000,-1038.8,-1503.0,-737.52,-1157.6
1774.000000000,83.190,1940.4,1992.4,1996.5,295.48,4462.6,967.00,11.415,6538.3,2753.7,3374.2,2098.2,0.0000,-6013.5,-6613.0,-946.96,-1808.3,-1241.3,-14814.,-90.793,-18547.,-5975.9,-3837.6,-2117.6,63.120,2248.6,2050.4,2108.6,325.83,4839.6,1686.6,0.0000,7740.9,4449.7,4252.8,3658.0,0.0000,-334.20,-101.59,-101.60,-42.080,-108.25,-587.69,0.0000,-1038.8,-1502.9,-737.49,-1157.5
1775.000000000,82.990,1934.7,1985.4,1995.5,294.72,4462.2,967.00,11.415,6538.4,2753.5,3374.1,2098.3,0.0000,-6010.1,-6610.8,-948.83,-1807.6,-1246.6,-14813.,-90.767,-18549.,-5975.6,-3837.3,-2117.2,62.932,2241.9,2044.3,2107.7,324.96,4839.6,1686.6,0.0000,7740.9,4449.7,4252.8,3658.0,0.0000,-333.14,-101.26,-101.50,-41.955,-108.42,-587.69,0.0000,-1038.8,-1502.9,-737.47,-1157.4
1776.000000000,82.793,1928.9,1979.4,1994.5,293.91,4462.2,967.00,11.415,6538.6,2753.1,3374.2,2098.4,0.0000,-6006.8,-6608.6,-950.64,-1807.0,-1251.7,-14813.,-90.740,-18551.,-5975.2,-3837.1,-2116.8,62.737,2235.0,2037.9,2106.9,324.05,4839.5,1686.6,0.0000,7740.9,4449.7,4252.8,3658.0,0.0000,-332.04,-100.91,-101.39,-41.825,-108.59,-587.69,0.0000,-1038.8,-1502.8,-737.44,-1157.3
1777.000000000,82.598,1923.0,1973.6,1993.6,293.26,4461.9,967.00,11.415,6560.1,2753.1,3374.1,2098.4,0.0000,-6003.3,-6606.4,-952.41,-1806.3,-1256.8,-14813.,-90.714,-18552.,-5974.9,-3836.9,-2116.4,62.611,2230.5,2033.8,2106.3,323.46,4839.4,1686.6,0.0000,7740.9,4449.7,4252.8,3658.0,0.0000,-331.30,-100.68,-101.33,-41.741,-108.76,-587.69,0.0000,-1038.8,-1502.8,-737.42,-1157.2
1778.000000000,82.442,1918.0,1968.5,1992.8,292.63,4461.5,966.99,10.128,6566.7,2752.8,3374.1,2098.5,0.0000,-5999.9,-6604.4,-954.13,-1805.6,-1261.7,-14813.,-90.687,-18554.,-5974.5,-3836.6,-2116.0,62.401,2223.0,2027.0,2105.4,322.48,4839.4,1686.6,0.0000,7740.9,4449.7,4252.8,3658.0,0.0000,-330.12,-100.31,-101.21,-41.601,-108.93,-587.69,0.0000,-1038.8,-1502.7,-737.39,-1157.1
1779.000000000,82.217,1914.7,1962.7,1991.9,291.83,4461.1,966.99,9.2206,6570.0,2752.8,3374.1,2098.6,0.0000,-5996.3,-6602.4,-955.81,-1804.9,-1266.5,-14812.,-90.661,-18555.,-5974.1,-3836.4,-2115.6,62.224,2216.7,2021.3,2104.6,321.65,4839.3,1686.6,0.0000,7740.9,4449.7,4252.8,3658.0,0.0000,-329.11,-99.999,-101.11,-41.483,-109.10,-587.69,0.0000,-1038.8,-1502.7,-737.37,-1157.0
1780.000000000,82.025,1909.0,1956.6,1991.1,291.03,4460.7,966.99,9.1976,6569.7,2752.8,3374.1,2098.6,0.0000,-5992.8,-6600.3,-957.45,-1804.2,-1271.2,-14812.,-90.634,-18557.,-5973.8,-3836.2,-2115.2,62.011,2209.1,2014.3,2103.6,320.66,4839.2,1686.6,0.0000,7740.9,4449.7,4252.8,3658.0,0.0000,-327.91,-99.625,-100.99,-41.340,-109.26,-587.69,0.0000,-1038.9,-1502.6,-737.35,-1156.9
1781.000000000,81.835,1903.1,1950.6,1990.3,290.20,4460.4,966.99,9.1976,6569.6,2752.9,3374.1,2098.7,0.0000,-5989.1,-6598.2,-959.03,-1803.5,-1275.8,-14812.,-90.608,-18558.,-5973.4,-3835.9,-2114.8,61.802,2201.7,2007.6,2102.7,319.68,4839.2,1686.6,0.0000,7740.9,4449.7,4252.8,3658.0,0.0000,-326.73,-99.259,-100.87,-41.201,-109.42,-587.69,0.0000,-1038.9,-1502.6,-737.32,-1156.8
1782.000000000,81.608,1896.8,1944.5,1994.0,289.43,4460.0,966.99,9.1976,6569.5,2753.0,3374.3,2098.7,0.0000,-5985.4,-6596.1,-960.58,-1802.8,-1280.4,-14812.,-90.581,-18559.,-5973.1,-3835.7,-2114.4,61.599,2194.4,2001.0,2101.8,318.74,4839.1,1686.6,0.0000,7740.9,4449.7,4252.8,3658.0,0.0000,-325.58,-98.903,-100.75,-41.066,-109.58,-587.69,0.0000,-1038.9,-1502.5,-737.30,-1156.7
1783.000000000,81.566,1890.7,1938.3,1999.0,288.59,4459.6,966.99,9.1976,6569.5,2753.0,3374.3,2098.8,0.0000,-5981.5,-6593.9,-962.09,-1802.1,-1284.8,-14811.,-90.555,-18560.,-5972.7,-3835.5,-2114.0,61.395,2187.2,1994.3,2100.9,317.78,4839.0,1686.6,0.0000,7740.9,4449.7,4252.8,3658.0,0.0000,-324.42,-98.543,-100.63,-40.930,-109.73,-587.69,0.0000,-1038.9,-1502.5,-737.27,-1156.6
1784.000000000,81.390,1884.9,1932.1,1998.2,287.87,4459.3,966.99,9.1976,6569.4,2753.1,3374.3,2098.9,0.0000,-5977.7,-6591.7,-963.56,-1801.4,-1289.2,-14811.,-90.528,-18561.,-5972.4,-3835.3,-2113.6,61.225,2181.1,1988.8,2100.1,316.99,4839.0,1686.6,0.0000,7740.9,4449.7,4252.8,3658.0,0.0000,-323.44,-98.239,-100.53,-40.817,-109.89,-587.69,0.0000,-1038.9,-1502.4,-737.25,-1156.5
1785.000000000,81.200,1879.3,1926.5,1997.2,287.17,4458.9,966.99,9.1976,6569.3,2753.1,3374.2,2099.0,0.0000,-5973.7,-6589.5,-965.00,-1800.7,-1293.4,-14811.,-90.502,-18562.,-5972.0,-3835.1,-2113.2,61.073,2175.7,1983.9,2099.4,316.28,4838.9,1686.6,0.0000,7740.9,4449.7,4252.8,3658.0,0.0000,-322.55,-97.963,-100.45,-40.715,-110.04,-587.69,0.0000,-1038.9,-1502.4,-737.23,-1156.4
1786.000000000,81.026,1874.2,1921.2,1996.5,286.43,4458.6,967.00,8.3418,6569.2,2753.2,3374.2,2099.1,0.0000,-5969.8,-6587.3,-966.40,-1800.0,-1297.6,-14811.,-90.475,-18563.,-5971.7,-3834.8,-2112.8,60.912,2170.0,1978.7,2098.7,315.53,4838.9,1686.6,0.0000,7740.9,4449.7,4252.8,3658.0,0.0000,-321.62,-97.674,-100.36,-40.608,-110.19,-587.69,0.0000,-1039.0,-1502.3,-737.20,-1156.3
1787.000000000,80.714,1868.9,1915.8,2000.1,285.76,4458.2,967.00,7.0151,6569.1,2753.2,3374.1,2099.1,0.0000,-5965.8,-6585.0,-967.77,-1799.2,-1301.8,-14810.,-90.449,-18564.,-5971.3,-3834.6,-2112.4,60.739,2163.8,1973.0,2097.9,314.72,4838.8,1686.6,0.0000,7740.9,4449.7,4252.8,3658.0,0.0000,-320.63,-97.365,-100.26,-40.493,-110.34,-587.69,0.0000,-1039.0,-1502.3,-737.18,-1156.2
1788.000000000,80.496,1863.8,1910.5,2005.4,285.10,4457.8,967.00,7.0153,6569.3,2753.3,3374.1,2099.2,0.0000,-5961.8,-6582.7,-969.11,-1798.5,-1305.8,-14810.,-90.422,-18565.,-5971.0,-3834.4,-2112.0,60.587,2158.4,1968.1,2097.3,314.01,4838.8,1686.6,0.0000,7740.9,4449.7,4252.8,3658.0,0.0000,-319.74,-97.089,-100.18,-40.391,-110.48,-587.69,0.0000,-1039.0,-1502.2,-737.16,-1156.1
1789.000000000,80.337,1858.7,1905.4,2004.4,284.48,4457.1,967.00,6.9968,6569.3,2753.3,3374.1,2099.3,0.0000,-5957.8,-6580.5,-970.41,-1797.8,-1309.8,-14810.,-90.396,-18566.,-5970.6,-3834.2,-2111.6,60.429,2152.7,1962.9,2092.9,313.21,4829.3,1686.6,0.0000,7735.1,4449.7,4252.8,3658.0,0.0000,-318.82,-96.804,-99.968,-40.286,-110.40,-587.69,0.0000,-1039.0,-1502.2,-737.13,-1156.0
1790.000000000,80.177,1853.7,1900.9,2002.5,283.80,4456.7,967.00,6.6721,6568.4,2753.3,3374.1,2099.3,0.0000,-5953.7,-6578.3,-971.64,-1797.1,-1313.6,-14810.,-90.369,-18567.,-5970.3,-3834.0,-2111.2,60.264,2146.9,1957.6,2086.1,312.34,4813.3,1686.6,0.0000,7725.5,4449.7,4252.8,3658.0,0.0000,-317.86,-96.509,-99.673,-40.176,-110.17,-587.69,0.0000,-1039.0,-1502.1,-737.11,-1155.9
1791.000000000,79.950,1848.8,1895.9,1999.2,283.06,4459.3,966.99,4.7983,6566.8,2753.4,3374.1,2099.4,0.0000,-5949.6,-6576.2,-972.81,-1796.3,-1317.2,-14809.,-90.342,-18568.,-5969.9,-3833.8,-2110.7,60.098,2141.0,1952.2,2079.1,311.46,4797.0,1686.6,0.0000,7715.6,4449.7,4252.8,3658.0,0.0000,-316.90,-96.212,-99.372,-40.066,-109.92,-587.69,0.0000,-1039.0,-1502.1,-737.09,-1155.8
1792.000000000,79.692,1844.0,1891.2,1994.4,282.31,4451.9,966.97,4.7986,6564.6,2753.5,3374.1,2099.5,0.0000,-5945.6,-6574.0,-973.89,-1795.6,-1320.7,-14809.,-90.316,-18569.,-5969.6,-3833.6,-2110.3,59.934,2135.1,1946.9,2072.0,310.58,4780.4,1686.6,0.0000,7705.5,4449.7,4252.8,3658.0,0.0000,-315.95,-95.918,-99.068,-39.956,-109.67,-587.69,0.0000,-1039.1,-1502.0,-737.07,-1155.7
1793.000000000,79.404,1839.2,1886.1,1988.9,281.53,4443.3,966.97,4.7990,6561.6,2753.5,3374.1,2099.6,0.0000,-5941.4,-6571.8,-974.88,-1794.9,-1324.0,-14809.,-90.289,-18569.,-5969.2,-3833.3,-2109.9,59.768,2129.2,1941.5,2064.7,309.70,4763.5,1686.6,0.0000,7695.3,4449.7,4252.8,3658.0,0.0000,-314.99,-95.621,-98.757,-39.846,-109.40,-587.69,0.0000,-1039.1,-1502.0,-737.04,-1155.6
1794.000000000,79.238,1834.8,1880.5,1982.8,280.75,4433.7,966.97,4.8033,6557.6,2753.6,3374.3,2099.6,0.0000,-5937.3,-6569.6,-975.78,-1794.1,-1327.2,-14808.,-90.263,-18570.,-5968.9,-3833.1,-2109.5,59.610,2123.6,1936.3,2057.6,308.85,4746.7,1686.6,0.0000,7685.1,4449.7,4252.8,3658.0,0.0000,-314.07,-95.336,-98.452,-39.740,-109.12,-587.69,0.0000,-1039.1,-1501.9,-737.02,-1155.5
1795.000000000,79.074,1830.2,1875.1,1976.4,280.01,4422.8,966.97,4.8037,6551.9,2753.7,3374.2,2099.7,0.0000,-5933.1,-6567.5,-976.59,-1793.4,-1330.2,-14808.,-90.236,-18571.,-5968.5,-3832.9,-2109.1,59.463,2118.3,1931.6,2050.6,308.06,4730.3,1686.6,0.0000,7675.1,4449.7,4252.8,3658.0,0.0000,-313.21,-95.069,-98.158,-39.642,-108.85,-587.69,0.0000,-1039.1,-1501.9,-737.00,-1155.4
1796.000000000,79.022,1825.8,1870.1,1970.1,279.29,4410.4,966.97,4.8172,6544.9,2753.7,3374.1,2099.6,0.0000,-5928.9,-6565.3,-977.34,-1792.7,-1333.1,-14808.,-90.209,-18571.,-5968.2,-3832.7,-2108.7,59.309,2112.8,1926.6,2043.4,307.22,4713.2,1686.6,0.0000,7664.8,4449.7,4252.8,3658.0,0.0000,-312.30,-94.790,-97.850,-39.539,-108.56,-587.69,0.0000,-1039.1,-1501.8,-736.97,-1155.3
1797.000000000,78.969,1821.0,1865.5,1963.7,278.56,4397.2,966.97,4.8200,6544.9,2753.4,3374.0,2099.6,0.0000,-5924.7,-6563.1,-978.01,-1791.9,-1335.8,-14807.,-90.183,-18572.,-5967.9,-3832.5,-2108.3,59.146,2107.0,1921.3,2035.9,306.35,4695.6,1686.6,0.0000,7654.1,4449.7,4252.8,3658.0,0.0000,-311.36,-94.498,-97.529,-39.431,-108.26,-587.69,0.0000,-1039.1,-1501.7,-736.95,-1155.2
1798.000000000,78.595,1816.1,1860.6,1957.0,277.81,4383.4,966.98,4.8203,6539.4,2753.5,3374.1,2099.7,0.0000,-5920.4,-6560.9,-978.61,-1791.2,-1338.4,-14807.,-90.156,-18572.,-5967.5,-3832.3,-2107.9,58.986,2101.4,1916.1,2028.4,305.49,4677.9,1686.6,0.0000,7643.3,4449.7,4252.8,3658.0,0.0000,-310.43,-94.211,-97.208,-39.324,-107.94,-587.69,0.0000,-1039.2,-1501.7,-736.93,-1155.1
1799.000000000,78.438,1811.1,1854.9,1950.2,277.06,4369.2,966.98,4.5017,6531.1,2753.5,3374.1,2099.8,0.0000,-5916.1,-6558.7,-979.15,-1790.4,-1341.0,-14807.,-90.130,-18573.,-5967.2,-3832.1,-2107.5,58.823,2095.5,1910.8,2020.7,304.60,4659.8,1686.6,0.0000,7632.4,4449.7,4252.8,3658.0,0.0000,-309.47,-93.918,-96.879,-39.215,-107.61,-587.69,0.0000,-1039.2,-1501.6,-736.91,-1155.0
1800.000000000,78.298,1806.4,1850.1,1951.3,276.32,4354.5,966.98,2.6054,6522.7,2753.6,3374.1,2099.8,0.0000,-5911.8,-6556.5,-979.62,-1789.7,-1343.4,-14806.,-90.103,-18573.,-5966.8,-3831.9,-2107.1,58.668,2090.0,1905.7,2013.2,303.76,4642.0,1686.6,0.0000,7621.6,4449.7,4252.8,3658.0,0.0000,-308.57,-93.638,-96.559,-39.112,-107.29,-587.69,0.0000,-1039.2,-1501.6,-736.88,-1154.9
1801.000000000,78.171,1803.1,1846.4,1946.8,275.78,4340.2,966.98,2.6059,6514.2,2753.5,3374.1,2099.8,0.0000,-5907.5,-6554.4,-980.07,-1789.0,-1345.6,-14806.,-90.077,-18574.,-5966.5,-3831.7,-2106.7,59.090,2096.0,1911.2,2012.1,304.62,4637.3,1686.6,0.0000,7618.6,4449.7,4252.8,3658.0,0.0000,-309.32,-93.870,-96.612,-39.220,-107.27,-587.69,0.0000,-1039.2,-1501.5,-736.86,-1154.8
1802.000000000,78.147,1808.2,1850.1,1941.6,276.71,4329.4,966.96,2.6065,6506.5,2753.3,3374.2,2099.9,0.0000,-5903.9,-6552.8,-980.59,-1788.3,-1347.9,-14806.,-90.053,-18574.,-5966.1,-3831.5,-2106.3,67.618,2152.6,1962.9,2031.8,313.13,4669.5,1686.6,5.5953,7639.0,4451.3,4254.1,3659.3,0.0000,-316.58,-96.209,-97.932,-40.160,-108.08,-587.69,-0.25547,-1039.2,-1501.5,-736.85,-1154.8
1803.000000000,78.732,1826.1,1865.3,1940.5,279.66,4325.1,966.90,2.6070,6500.5,2753.3,3374.2,2100.0,0.0000,-5901.5,-6551.9,-981.18,-1787.8,-1350.3,-14805.,-90.029,-18574.,-5965.8,-3831.3,-2105.9,106.69,2245.2,2023.8,2045.9,321.24,4676.8,1686.6,66.363,7648.8,4457.7,4262.3,3667.1,0.0000,-319.81,-98.042,-98.325,-40.597,-108.17,-587.69,-3.0300,-1039.4,-1501.4,-736.86,-1154.8
1804.000000000,79.300,1843.7,1881.9,1942.4,281.54,4321.8,966.90,2.6076,6495.3,2753.4,3374.1,2100.1,0.0000,-5900.2,-6551.9,-981.84,-1787.4,-1352.9,-14805.,-90.005,-18575.,-5965.5,-3831.1,-2105.5,61.360,2185.9,1993.2,2029.3,316.48,4653.4,1686.6,0.0000,7628.0,4449.7,4252.9,3658.1,0.0000,-322.43,-97.860,-98.513,-40.907,-107.90,-587.69,0.0000,-1039.2,-1501.4,-736.79,-1154.6
1805.000000000,79.813,1856.8,1894.6,1943.7,283.96,4315.2,966.90,2.6082,6489.6,2753.4,3374.1,2100.2,0.0000,-5899.5,-6552.1,-982.51,-1787.1,-1355.2,-14805.,-89.980,-18575.,-5965.1,-3830.9,-2105.1,61.486,2190.4,1997.3,2023.6,316.95,4637.1,1686.6,0.0000,7618.1,4449.7,4252.9,3658.1,0.0000,-323.03,-98.054,-98.397,-40.991,-107.60,-587.69,0.0000,-1039.3,-1501.3,-736.77,-1154.5
1806.000000000,80.412,1863.8,1902.2,1942.9,285.31,4316.0,966.90,2.6087,6484.2,2753.5,3374.1,2100.3,0.0000,-5899.0,-6552.3,-983.22,-1786.8,-1357.4,-14804.,-89.954,-18575.,-5964.8,-3830.7,-2104.7,61.498,2190.8,1997.7,2022.1,316.98,4633.3,1686.6,0.0000,7615.7,4449.7,4252.9,3658.1,0.0000,-323.05,-98.068,-98.363,-40.999,-107.59,-587.69,0.0000,-1039.3,-1501.3,-736.75,-1154.4
1807.000000000,80.645,1866.8,1906.3,1940.7,285.94,4308.4,966.90,2.6093,6481.1,2753.5,3374.3,2100.4,0.0000,-5898.4,-6552.4,-983.89,-1786.4,-1359.6,-14804.,-89.928,-18575.,-5964.4,-3830.5,-2104.3,61.452,2189.2,1996.2,2020.6,316.72,4629.9,1686.6,0.0000,7613.7,4449.7,4252.8,3658.0,0.0000,-322.76,-97.990,-98.297,-40.968,-107.60,-587.69,0.0000,-1039.3,-1501.2,-736.73,-1154.3
1808.000000000,80.768,1867.9,1907.2,1938.1,286.07,4305.2,966.90,2.6098,6480.8,2753.6,3374.3,2100.5,0.0000,-5897.7,-6552.4,-984.48,-1786.0,-1361.6,-14803.,-89.902,-18576.,-5964.1,-3830.3,-2103.8,61.381,2186.7,1993.9,2019.1,316.34,4626.6,1686.6,0.0000,7611.7,4449.7,4252.8,3658.0,0.0000,-322.35,-97.872,-98.215,-40.921,-107.60,-587.69,0.0000,-1039.3,-1501.2,-736.71,-1154.2
1809.000000000,80.756,1867.6,1907.7,1935.9,285.89,4303.5,966.90,2.6103,6479.1,2753.6,3374.3,2100.5,0.0000,-5896.8,-6552.1,-985.02,-1785.6,-1363.7,-14803.,-89.876,-18576.,-5963.7,-3830.0,-2103.4,61.288,2183.4,1990.9,2017.4,315.88,4623.3,1686.6,0.0000,7609.7,4449.7,4252.8,3658.0,0.0000,-321.81,-97.718,-98.117,-40.859,-107.60,-587.69,0.0000,-1039.3,-1501.1,-736.68,-1154.1
1810.000000000,80.695,1866.2,1907.6,1934.4,285.56,4300.6,966.90,2.6108,6475.3,2753.7,3374.3,2100.5,0.0000,-5895.8,-6551.8,-985.54,-1785.2,-1365.7,-14803.,-89.850,-18576.,-5963.4,-3829.8,-2103.0,61.181,2179.6,1987.4,2015.6,315.35,4619.9,1686.6,0.0000,7607.7,4449.7,4252.8,3658.0,0.0000,-321.21,-97.540,-98.010,-40.788,-107.60,-587.69,0.0000,-1039.3,-1501.1,-736.66,-1154.0
1811.000000000,80.608,1865.4,1907.0,1933.3,285.21,4302.4,966.90,2.6114,6470.6,2753.8,3374.3,2100.7,0.0000,-5894.7,-6551.4,-986.05,-1784.7,-1367.6,-14802.,-89.823,-18576.,-5963.0,-3829.6,-2102.6,61.100,2176.7,1984.8,2014.1,314.95,4616.9,1686.6,0.0000,7605.8,4449.7,4252.8,3658.0,0.0000,-320.74,-97.403,-97.924,-40.734,-107.61,-587.69,0.0000,-1039.3,-1501.0,-736.64,-1153.9
1812.000000000,80.432,1864.9,1906.5,1932.4,285.05,4296.8,966.91,2.6119,6466.6,2753.8,3374.4,2100.8,0.0000,-5893.5,-6550.9,-986.56,-1784.2,-1369.5,-14802.,-89.798,-18576.,-5962.7,-3829.4,-2102.2,71.738,2243.8,2006.3,2035.6,317.96,4629.2,1686.6,48.381,7623.6,4459.1,4264.8,3669.0,0.0000,-321.80,-98.028,-98.054,-40.875,-107.74,-587.69,-2.2090,-1039.6,-1501.0,-736.67,-1153.9
1813.000000000,80.407,1866.6,1907.0,1931.4,285.20,4293.3,966.91,2.6124,6463.9,2753.9,3374.4,2100.8,0.0000,-5892.3,-6550.6,-987.06,-1783.8,-1371.4,-14801.,-89.772,-18576.,-5962.3,-3829.2,-2101.8,61.215,2180.7,1988.5,2013.2,315.46,4613.3,1686.6,0.0000,7603.6,4449.7,4252.8,3658.0,0.0000,-321.25,-97.568,-97.966,-40.810,-107.68,-587.69,0.0000,-1039.4,-1500.9,-736.59,-1153.7
1814.000000000,80.355,1867.4,1907.0,1930.8,284.94,4290.5,966.91,2.6129,6461.7,2753.9,3374.6,2100.9,0.0000,-5891.0,-6550.2,-987.57,-1783.4,-1373.3,-14801.,-89.747,-18577.,-5962.0,-3829.0,-2101.4,61.174,2179.3,1987.2,2011.9,315.25,4610.5,1686.6,0.0000,7601.9,4449.7,4252.8,3658.0,0.0000,-320.99,-97.495,-97.909,-40.783,-107.69,-587.69,0.0000,-1039.4,-1500.9,-736.57,-1153.6
1815.000000000,80.064,1866.7,1906.2,1930.1,284.90,4287.0,966.91,2.6134,6459.3,2754.0,3374.7,2101.1,0.0000,-5889.6,-6549.8,-988.07,-1782.9,-1375.1,-14800.,-89.721,-18577.,-5961.6,-3828.8,-2101.0,61.061,2175.2,1983.5,2010.1,314.70,4607.0,1686.6,0.0000,7599.9,4449.7,4252.8,3658.0,0.0000,-320.35,-97.305,-97.796,-40.707,-107.68,-587.69,0.0000,-1039.4,-1500.8,-736.55,-1153.5
1816.000000000,80.044,1864.9,1904.5,1928.9,284.57,4282.9,966.92,2.6139,6457.0,2754.0,3374.7,2101.2,0.0000,-5888.1,-6549.3,-988.55,-1782.5,-1376.9,-14800.,-89.695,-18577.,-5961.3,-3828.6,-2100.6,60.925,2170.4,1979.1,2008.2,314.04,4603.5,1686.6,0.0000,7597.7,4449.7,4252.8,3658.0,0.0000,-319.59,-97.079,-97.666,-40.617,-107.67,-587.69,0.0000,-1039.4,-1500.8,-736.53,-1153.4
1817.000000000,79.934,1862.5,1902.3,1927.4,284.10,4278.9,966.92,2.6145,6454.8,2754.1,3375.0,2101.2,0.0000,-5886.4,-6548.8,-989.01,-1782.0,-1378.6,-14799.,-89.669,-18577.,-5960.9,-3828.4,-2100.2,60.772,2165.0,1974.1,2006.1,313.30,4599.8,1686.6,0.0000,7595.5,4449.7,4252.8,3658.0,0.0000,-318.74,-96.822,-97.523,-40.514,-107.66,-587.69,0.0000,-1039.4,-1500.7,-736.51,-1153.3
1818.000000000,79.990,1859.2,1899.8,1925.7,283.54,4275.4,966.92,2.6150,6452.8,2753.8,3375.1,2101.2,0.0000,-5884.6,-6548.2,-989.45,-1781.5,-1380.4,-14799.,-89.643,-18577.,-5960.6,-3828.2,-2099.8,60.663,2161.1,1970.6,2005.2,312.79,4598.7,1686.6,0.0000,7594.9,4449.7,4252.8,3658.0,0.0000,-318.12,-96.638,-97.443,-40.442,-107.70,-587.69,0.0000,-1039.4,-1500.7,-736.48,-1153.2
1819.000000000,79.875,1856.2,1896.9,1924.2,283.04,4272.4,966.92,2.6155,6450.8,2753.8,3375.1,2101.3,0.0000,-5882.8,-6547.5,-989.87,-1781.0,-1382.1,-14798.,-89.617,-18577.,-5960.2,-3828.0,-2099.4,60.536,2156.5,1966.4,2004.4,312.19,4598.2,1686.6,0.0000,7594.6,4449.7,4252.8,3658.0,0.0000,-317.40,-96.421,-97.357,-40.357,-107.76,-587.69,0.0000,-1039.5,-1500.6,-736.46,-1153.1
1820.000000000,79.746,1853.1,1893.9,1923.0,282.49,4269.8,966.92,2.6160,6449.2,2753.9,3375.3,2101.4,0.0000,-5880.9,-6546.7,-990.29,-1780.5,-1383.8,-14798.,-89.590,-18577.,-5959.9,-3827.8,-2099.0,60.410,2152.1,1962.3,2003.7,311.60,4597.7,1686.6,0.0000,7594.3,4449.7,4252.8,3658.0,0.0000,-316.69,-96.206,-97.273,-40.273,-107.82,-587.69,0.0000,-1039.5,-1500.6,-736.44,-1153.0
1821.000000000,79.625,1849.9,1890.4,1922.1,281.99,4267.4,966.92,2.6165,6447.7,2753.9,3375.4,2101.5,0.0000,-5878.8,-6545.9,-990.70,-1780.0,-1385.5,-14798.,-89.564,-18577.,-5959.5,-3827.6,-2098.6,60.287,2147.7,1958.3,2003.0,311.02,4597.2,1686.6,0.0000,7594.1,4449.7,4252.8,3658.0,0.0000,-315.99,-95.996,-97.191,-40.191,-107.88,-587.69,0.0000,-1039.5,-1500.5,-736.42,-1152.9
1822.000000000,79.547,1846.6,1886.7,1921.4,281.51,4265.4,966.92,2.6169,6446.0,2754.0,3375.6,2101.6,0.0000,-5876.7,-6545.0,-991.11,-1779.5,-1387.1,-14797.,-89.538,-18577.,-5959.2,-3827.4,-2098.2,60.189,2144.2,1955.2,2002.4,310.56,4596.8,1686.6,0.0000,7593.8,4449.7,4252.8,3658.0,0.0000,-315.42,-95.825,-97.126,-40.126,-107.94,-587.69,0.0000,-1039.5,-1500.5,-736.40,-1152.8
1823.000000000,79.432,1843.6,1883.4,1920.9,281.08,4263.5,966.92,2.6174,6444.4,2753.8,3375.6,2101.7,0.0000,-5874.4,-6544.0,-991.51,-1778.9,-1388.8,-14797.,-89.512,-18577.,-5958.9,-3827.2,-2097.8,60.099,2141.0,1952.2,2001.8,310.14,4596.4,1686.6,0.0000,7593.6,4449.7,4252.8,3658.0,0.0000,-314.89,-95.666,-97.066,-40.066,-107.99,-587.69,0.0000,-1039.5,-1500.4,-736.37,-1152.7
1824.000000000,79.328,1840.7,1880.5,1920.4,280.62,4261.8,966.92,2.6179,6443.0,2753.6,3375.8,2101.8,0.0000,-5872.1,-6543.0,-991.91,-1778.4,-1390.5,-14796.,-89.486,-18577.,-5958.5,-3827.0,-2097.4,59.979,2136.7,1948.3,2001.1,309.58,4595.9,1686.6,0.0000,7593.3,4449.7,4252.8,3658.0,0.0000,-314.21,-95.458,-96.985,-39.986,-108.05,-587.69,0.0000,-1039.5,-1500.4,-736.35,-1152.6
1825.000000000,79.215,1837.4,1877.3,1920.0,280.15,4260.5,966.93,2.6184,6441.9,2753.5,3375.7,2101.9,0.0000,-5869.7,-6542.0,-992.31,-1777.9,-1392.2,-14796.,-89.460,-18577.,-5958.1,-3826.8,-2097.0,59.851,2132.2,1944.2,2000.4,308.98,4595.4,1686.6,0.0000,7593.0,4449.7,4252.8,3658.0,0.0000,-313.48,-95.237,-96.899,-39.901,-108.11,-587.69,0.0000,-1039.5,-1500.3,-736.33,-1152.5
1826.000000000,79.098,1833.8,1873.8,1919.5,279.68,4259.4,966.93,2.6189,6441.0,2753.5,3375.8,2102.0,0.0000,-5867.2,-6540.9,-992.70,-1777.3,-1393.8,-14795.,-89.434,-18577.,-5957.8,-3826.6,-2096.6,59.713,2127.2,1939.7,1999.6,308.33,4594.9,1686.6,0.0000,7592.7,4449.7,4252.8,3658.0,0.0000,-312.69,-94.999,-96.806,-39.809,-108.16,-587.69,0.0000,-1039.5,-1500.3,-736.31,-1152.4
1827.000000000,78.975,1830.2,1870.8,1918.9,279.17,4258.4,966.93,2.6194,6440.2,2753.6,3375.9,2102.1,0.0000,-5864.6,-6539.8,-993.08,-1776.8,-1395.4,-14795.,-89.408,-18577.,-5957.4,-3826.4,-2096.2,59.609,2123.5,1936.3,1999.0,307.84,4594.4,1686.6,0.0000,7592.5,4449.7,4252.8,3658.0,0.0000,-312.08,-94.814,-96.736,-39.739,-108.22,-587.69,0.0000,-1039.5,-1500.2,-736.29,-1152.3
1828.000000000,78.856,1827.0,1868.3,1918.2,278.73,4257.6,966.93,2.6198,6439.5,2753.7,3375.9,2102.2,0.0000,-5862.1,-6538.6,-993.46,-1776.2,-1397.1,-14794.,-89.382,-18577.,-5957.1,-3826.2,-2095.8,59.540,2121.1,1934.1,1998.6,307.52,4594.2,1686.6,0.0000,7592.3,4449.7,4252.8,3658.0,0.0000,-311.66,-94.686,-96.692,-39.693,-108.27,-587.69,0.0000,-1039.6,-1500.1,-736.26,-1152.3
1829.000000000,78.757,1824.4,1866.0,1917.5,278.35,4256.6,966.93,2.6203,6439.0,2753.7,3375.8,2102.3,0.0000,-5859.6,-6537.4,-993.84,-1775.7,-1398.6,-14793.,-89.356,-18577.,-5956.7,-3826.0,-2095.4,59.451,2117.9,1931.2,1998.2,307.10,4594.1,1686.6,0.0000,7592.3,4449.7,4252.8,3658.0,0.0000,-311.13,-94.525,-96.637,-39.634,-108.34,-587.69,0.0000,-1039.6,-1500.1,-736.24,-1152.2
1830.000000000,78.658,1821.7,1863.3,1917.0,277.94,4255.8,966.93,2.6208,6438.5,2753.8,3375.7,2102.4,0.0000,-5857.0,-6536.2,-994.21,-1775.1,-1400.2,-14793.,-89.330,-18577.,-5956.4,-3825.8,-2095.0,59.335,2113.8,1927.4,1997.6,306.56,4594.0,1686.6,0.0000,7592.3,4449.7,4252.8,3658.0,0.0000,-310.46,-94.322,-96.565,-39.557,-108.40,-587.69,0.0000,-1039.6,-1500.0,-736.22,-1152.1
1831.000000000,78.554,1818.6,1860.3,1916.7,277.57,4255.3,966.93,2.6213,6438.0,2753.8,3375.7,2102.5,0.0000,-5854.5,-6534.9,-994.57,-1774.6,-1401.8,-14792.,-89.304,-18577.,-5956.0,-3825.6,-2094.5,59.210,2109.3,1923.4,1997.0,305.98,4594.0,1686.6,0.0000,7592.3,4449.7,4252.8,3658.0,0.0000,-309.74,-94.103,-96.486,-39.473,-108.46,-587.69,0.0000,-1039.6,-1500.0,-736.20,-1152.0
1832.000000000,78.447,1815.0,1857.2,1916.2,277.08,4254.7,966.93,2.6218,6437.4,2753.9,3375.8,2102.5,0.0000,-5851.8,-6533.6,-994.93,-1774.0,-1403.4,-14792.,-89.278,-18577.,-5955.6,-3825.4,-2094.1,59.075,2104.5,1919.0,1996.4,305.34,4593.9,1686.6,0.0000,7592.2,4449.7,4252.8,3658.0,0.0000,-308.97,-93.867,-96.400,-39.383,-108.52,-587.69,0.0000,-1039.6,-1499.9,-736.18,-1151.9
1833.000000000,78.330,1811.1,1853.9,1915.8,276.57,4254.1,966.93,2.6222,6437.0,2753.9,3375.9,2102.6,0.0000,-5849.1,-6532.2,-995.28,-1773.4,-1404.9,-14791.,-89.252,-18577.,-5955.3,-3825.2,-2093.7,58.941,2099.8,1914.6,1995.8,304.72,4593.8,1686.6,0.0000,7592.2,4449.7,4252.8,3658.0,0.0000,-308.20,-93.634,-96.315,-39.294,-108.58,-587.69,0.0000,-1039.6,-1499.9,-736.15,-1151.8
1834.000000000,78.194,1806.8,1850.2,1915.3,276.10,4260.2,966.93,2.6227,6436.8,2753.7,3375.9,2102.7,0.0000,-5846.4,-6530.8,-995.62,-1772.8,-1406.5,-14791.,-89.226,-18577.,-5954.9,-3825.0,-2093.3,58.805,2094.9,1910.2,1995.2,304.08,4593.7,1686.6,0.0000,7592.2,4449.7,4252.8,3658.0,0.0000,-307.42,-93.396,-96.229,-39.203,-108.64,-587.69,0.0000,-1039.6,-1499.8,-736.13,-1151.7
1835.000000000,77.871,1802.9,1846.2,1914.7,275.55,4263.3,966.93,2.6231,6436.6,2753.7,3375.8,2102.8,0.0000,-5843.5,-6529.4,-995.96,-1772.3,-1408.0,-14790.,-89.200,-18577.,-5954.6,-3824.8,-2092.9,58.665,2089.9,1905.7,1994.6,303.43,4593.6,1686.6,0.0000,7592.2,4449.7,4252.8,3658.0,0.0000,-306.62,-93.152,-96.140,-39.110,-108.70,-587.69,0.0000,-1039.6,-1499.8,-736.11,-1151.6
1836.000000000,77.739,1799.1,1842.3,1914.1,275.00,4262.9,966.90,2.6236,6436.2,2753.8,3375.7,2102.9,0.0000,-5840.6,-6527.9,-996.29,-1771.7,-1409.5,-14790.,-89.174,-18577.,-5954.2,-3824.6,-2092.5,58.523,2084.9,1901.0,1993.9,302.77,4593.6,1686.6,0.0000,7592.2,4449.7,4252.8,3658.0,0.0000,-305.81,-92.904,-96.049,-39.015,-108.76,-587.69,0.0000,-1039.6,-1499.7,-736.09,-1151.5
1837.000000000,77.599,1795.3,1838.4,1913.5,274.41,4262.5,966.89,2.6241,6435.9,2753.8,3375.7,2103.0,0.0000,-5837.6,-6526.4,-996.61,-1771.1,-1411.0,-14789.,-89.148,-18577.,-5953.9,-3824.4,-2092.1,58.377,2079.7,1896.3,1993.3,302.09,4593.5,1686.6,0.0000,7592.2,4449.7,4252.8,3658.0,0.0000,-304.97,-92.649,-95.957,-38.918,-108.82,-587.69,0.0000,-1039.7,-1499.7,-736.07,-1151.4
1838.000000000,77.456,1791.2,1834.0,1913.0,273.83,4262.1,966.89,2.6245,6435.6,2753.7,3375.5,2103.2,0.0000,-5834.5,-6524.9,-996.93,-1770.5,-1412.5,-14789.,-89.122,-18577.,-5953.5,-3824.2,-2091.7,58.254,2075.3,1892.3,1992.7,301.52,4593.4,1686.6,0.0000,7592.2,4449.7,4252.8,3658.0,0.0000,-304.26,-92.431,-95.879,-38.836,-108.87,-587.69,0.0000,-1039.7,-1499.6,-736.04,-1151.3
1839.000000000,77.102,1787.4,1829.8,1912.4,273.30,4261.7,966.89,2.6250,6435.5,2753.6,3375.2,2103.3,0.0000,-5831.3,-6523.3,-997.23,-1769.8,-1414.0,-14788.,-89.096,-18577.,-5953.2,-3824.0,-2091.3,58.134,2071.0,1888.4,1992.2,300.95,4593.4,1686.6,0.0000,7592.2,4449.7,4252.8,3658.0,0.0000,-303.56,-92.216,-95.804,-38.756,-108.93,-587.69,0.0000,-1039.7,-1499.6,-736.02,-1151.2
1840.000000000,76.669,1783.8,1825.9,1911.8,272.78,4261.3,966.90,2.6258,6435.3,2753.6,3375.2,2103.3,0.0000,-5828.1,-6521.7,-997.54,-1769.2,-1415.5,-14788.,-89.069,-18577.,-5952.8,-3823.8,-2090.9,58.016,2066.8,1884.6,1991.6,300.40,4593.4,1686.6,0.0000,7592.2,4449.7,4252.8,3658.0,0.0000,-302.87,-92.005,-95.730,-38.677,-108.99,-587.69,0.0000,-1039.7,-1499.5,-736.00,-1151.1
1841.000000000,76.524,1780.2,1822.1,1911.2,272.29,4261.0,966.87,2.6288,6435.0,2753.7,3375.1,2103.3,0.0000,-5824.9,-6520.1,-997.84,-1768.6,-1416.9,-14787.,-89.043,-18577.,-5952.5,-3823.6,-2090.5,57.893,2062.4,1880.6,1991.1,299.83,4593.3,1686.6,0.0000,7592.2,4449.7,4252.8,3658.0,0.0000,-302.15,-91.786,-95.652,-38.596,-109.04,-587.69,0.0000,-1039.7,-1499.5,-735.98,-1151.0
1842.000000000,76.402,1776.7,1818.5,1910.6,271.82,4260.7,966.85,2.6040,6434.9,2753.5,3374.9,2103.4,0.0000,-5821.6,-6518.6,-998.13,-1768.0,-1418.4,-14786.,-89.018,-18577.,-5952.1,-3823.4,-2090.1,57.795,2058.9,1877.4,1990.6,299.37,4593.3,1686.6,0.0000,7592.1,4449.7,4252.8,3658.0,0.0000,-301.56,-91.607,-95.591,-38.530,-109.10,-587.69,0.0000,-1039.7,-1499.4,-735.96,-1150.9
1843.000000000,76.331,1773.6,1815.1,1910.1,271.40,4260.4,966.85,2.5964,6434.7,2753.5,3374.9,2103.7,0.0000,-5818.3,-6517.0,-998.42,-1767.4,-1419.8,-14786.,-88.992,-18577.,-5951.8,-3823.1,-2089.7,57.706,2055.7,1874.5,1990.2,298.96,4593.3,1686.6,0.0000,7592.1,4449.7,4252.8,3658.0,0.0000,-301.02,-91.441,-95.536,-38.471,-109.15,-587.69,0.0000,-1039.7,-1499.4,-735.93,-1150.8
1844.000000000,76.286,1770.8,1811.9,1909.5,270.98,4260.2,966.85,2.5968,6434.6,2753.5,3374.7,2103.8,0.0000,-5815.1,-6515.4,-998.70,-1766.8,-1421.2,-14785.,-88.966,-18577.,-5951.4,-3822.9,-2089.3,57.608,2052.3,1871.3,1989.8,298.50,4593.2,1686.6,0.0000,7592.1,4449.7,4252.8,3658.0,0.0000,-300.43,-91.262,-95.475,-38.406,-109.21,-587.69,0.0000,-1039.7,-1499.3,-735.91,-1150.7
1845.000000000,76.182,1767.8,1808.8,1909.0,270.58,4259.9,966.85,2.5973,6434.4,2753.6,3374.7,2103.8,0.0000,-5811.8,-6513.8,-998.98,-1766.1,-1422.6,-14785.,-88.940,-18577.,-5951.1,-3822.7,-2088.9,57.521,2049.2,1868.5,1989.4,298.09,4593.2,1686.6,0.0000,7592.1,4449.7,4252.8,3658.0,0.0000,-299.90,-91.100,-95.422,-38.348,-109.26,-587.69,0.0000,-1039.7,-1499.3,-735.89,-1150.6
1846.000000000,75.893,1764.8,1805.3,1908.4,270.17,4259.3,966.85,2.5977,6434.2,2753.6,3374.7,2103.9,0.0000,-5808.5,-6512.2,-999.25,-1765.5,-1424.0,-14784.,-88.914,-18577.,-5950.7,-3822.5,-2088.5,57.409,2045.2,1864.8,1986.3,297.53,4586.5,1686.6,0.0000,7588.1,4449.7,4252.8,3658.0,0.0000,-299.24,-90.898,-95.266,-38.273,-109.15,-587.69,0.0000,-1039.7,-1499.2,-735.87,-1150.5
1847.000000000,75.712,1761.8,1801.9,1906.8,269.69,4256.5,966.85,2.5982,6433.5,2753.7,3374.8,2104.0,0.0000,-5805.2,-6510.7,-999.45,-1764.9,-1425.3,-14784.,-88.888,-18577.,-5950.4,-3822.3,-2088.1,57.263,2040.0,1860.1,1972.8,296.63,4553.0,1686.6,0.0000,7567.7,4449.7,4252.8,3658.0,0.0000,-298.40,-90.643,-94.749,-38.176,-108.39,-587.69,0.0000,-1039.8,-1499.2,-735.85,-1150.4
1848.000000000,75.591,1758.0,1798.1,1902.2,269.08,4248.2,966.85,2.5986,6431.3,2753.8,3375.0,2104.0,0.0000,-5801.8,-6509.1,-999.57,-1764.3,-1426.4,-14783.,-88.862,-18577.,-5950.0,-3822.1,-2087.7,57.124,2035.0,1855.6,1959.5,295.76,4520.1,1686.6,0.0000,7547.8,4449.7,4252.8,3658.0,0.0000,-297.60,-90.398,-94.242,-38.083,-107.63,-587.69,0.0000,-1039.8,-1499.1,-735.82,-1150.3
1849.000000000,75.472,1754.2,1794.1,1894.8,268.37,4235.0,966.85,2.5990,6427.4,2753.8,3375.0,2104.1,0.0000,-5798.3,-6507.4,-999.59,-1763.7,-1427.2,-14782.,-88.836,-18577.,-5949.7,-3821.9,-2087.3,57.008,2030.9,1851.8,1947.0,295.01,4488.8,1686.6,0.0000,7528.8,4449.7,4252.8,3658.0,0.0000,-296.91,-90.188,-93.770,-38.005,-106.91,-587.69,0.0000,-1039.8,-1499.0,-735.80,-1150.2
1850.000000000,75.319,1750.4,1790.4,1885.5,267.62,4227.0,966.85,2.5995,6422.2,2753.9,3375.1,2104.2,0.0000,-5794.8,-6505.8,-999.49,-1763.0,-1427.8,-14782.,-88.811,-18577.,-5949.4,-3821.7,-2086.9,56.889,2026.7,1848.0,1934.5,294.25,4457.6,1686.6,0.0000,7509.8,4449.7,4252.8,3658.0,0.0000,-296.21,-89.976,-93.298,-37.926,-106.19,-587.69,0.0000,-1039.8,-1499.0,-735.78,-1150.1
1851.000000000,75.091,1747.0,1786.7,1875.1,266.89,4212.5,966.85,2.5999,6415.6,2753.9,3375.0,2104.3,0.0000,-5791.3,-6504.1,-999.26,-1762.4,-1428.3,-14781.,-88.785,-18577.,-5949.0,-3821.4,-2086.5,56.769,2022.4,1844.1,1922.0,293.49,4426.5,1686.6,0.0000,7491.0,4449.7,4252.8,3658.0,0.0000,-295.51,-89.760,-92.823,-37.846,-105.46,-587.69,0.0000,-1039.8,-1498.9,-735.76,-1150.0
1852.000000000,74.973,1743.8,1783.3,1864.1,266.19,4194.1,966.85,2.6003,6406.7,2754.0,3375.0,2104.4,0.0000,-5787.8,-6502.5,-998.90,-1761.7,-1428.5,-14781.,-88.759,-18577.,-5948.7,-3821.2,-2086.1,56.652,2018.2,1840.3,1909.7,292.74,4395.8,1686.6,0.0000,7472.3,4449.7,4252.8,3658.0,0.0000,-294.81,-89.550,-92.355,-37.768,-104.74,-587.69,0.0000,-1039.8,-1498.9,-735.74,-1149.9
1853.000000000,74.727,1740.3,1779.6,1853.1,265.53,4172.6,966.85,2.6007,6394.4,2754.0,3375.0,2104.5,0.0000,-5784.2,-6500.8,-998.44,-1761.1,-1428.6,-14780.,-88.733,-18576.,-5948.3,-3821.0,-2085.7,56.511,2013.2,1835.7,1896.8,291.87,4363.9,1686.6,0.0000,7453.0,4449.7,4252.8,3658.0,0.0000,-294.00,-89.301,-91.855,-37.674,-103.98,-587.69,0.0000,-1039.8,-1498.8,-735.72,-1149.8
1854.000000000,74.498,1736.8,1775.7,1842.1,264.80,4148.1,966.85,2.6012,6380.2,2754.1,3375.0,2104.6,0.0000,-5780.6,-6499.1,-997.89,-1760.4,-1428.6,-14780.,-88.707,-18576.,-5948.0,-3820.8,-2085.3,56.385,2008.7,1831.6,1884.4,291.08,4333.1,1686.6,0.0000,7434.2,4449.7,4252.8,3658.0,0.0000,-293.26,-89.076,-91.377,-37.590,-103.25,-587.69,0.0000,-1039.8,-1498.8,-735.69,-1149.7
1855.000000000,74.373,1733.0,1771.7,1830.8,264.10,4123.1,966.86,2.6016,6365.4,2754.1,3375.1,2104.7,0.0000,-5777.0,-6497.5,-997.27,-1759.8,-1428.5,-14779.,-88.682,-18576.,-5947.6,-3820.6,-2084.9,56.259,2004.2,1827.5,1872.1,290.29,4302.5,1686.6,0.0000,7415.7,4449.7,4252.8,3658.0,0.0000,-292.52,-88.851,-90.902,-37.506,-102.51,-587.69,0.0000,-1039.8,-1498.7,-735.67,-1149.6
1856.000000000,74.324,1729.3,1768.0,1819.2,263.37,4098.1,966.86,2.6020,6350.4,2754.3,3375.3,2104.7,0.0000,-5773.3,-6495.8,-996.56,-1759.1,-1428.2,-14778.,-88.656,-18575.,-5947.3,-3820.4,-2084.5,56.136,1999.8,1823.5,1859.9,289.52,4272.3,1686.6,0.0000,7397.3,4449.7,4252.8,3658.0,0.0000,-291.80,-88.631,-90.433,-37.424,-101.78,-587.69,0.0000,-1039.8,-1498.7,-735.65,-1149.5
1857.000000000,74.168,1725.6,1764.2,1807.8,262.66,4073.2,966.86,2.6024,6335.6,2754.5,3375.4,2104.8,0.0000,-5769.6,-6494.1,-995.79,-1758.5,-1427.9,-14778.,-88.630,-18575.,-5946.9,-3820.2,-2084.1,56.013,1995.4,1819.5,1847.8,288.75,4242.3,1686.6,0.0000,7379.1,4449.7,4252.8,3658.0,0.0000,-291.08,-88.411,-89.966,-37.342,-101.06,-587.69,0.0000,-1039.8,-1498.6,-735.63,-1149.4
1858.000000000,73.971,1721.8,1760.3,1796.6,261.95,4048.0,966.86,2.6028,6320.5,2754.6,3375.5,2104.8,0.0000,-5765.8,-6492.4,-994.94,-1757.8,-1427.4,-14777.,-88.604,-18575.,-5946.6,-3819.9,-2083.7,55.874,1990.5,1815.0,1835.4,287.90,4211.6,1686.6,0.0000,7360.4,4449.7,4252.8,3658.0,0.0000,-290.27,-88.165,-89.478,-37.249,-100.31,-587.69,0.0000,-1039.9,-1498.6,-735.61,-1149.3
1859.000000000,73.840,1717.8,1756.2,1785.4,261.22,4022.1,966.86,2.6032,6305.1,2754.5,3375.6,2104.9,0.0000,-5762.1,-6490.7,-994.03,-1757.2,-1426.7,-14776.,-88.579,-18574.,-5946.2,-3819.7,-2083.3,55.743,1985.8,1810.7,1823.2,287.08,4181.4,1686.6,0.0000,7342.1,4449.7,4252.8,3658.0,0.0000,-289.50,-87.931,-89.002,-37.162,-99.567,-587.69,0.0000,-1039.9,-1498.5,-735.59,-1149.2
1860.000000000,73.708,1714.0,1752.3,1774.0,260.51,3996.1,966.86,2.6037,6289.8,2754.3,3375.7,2105.0,0.0000,-5758.3,-6488.9,-993.07,-1756.5,-1426.0,-14776.,-88.553,-18574.,-5945.9,-3819.5,-2082.9,55.636,1982.0,1807.3,1811.7,286.40,4152.8,1686.6,0.0000,7324.7,4449.7,4252.8,3658.0,0.0000,-288.87,-87.736,-88.562,-37.091,-98.862,-587.69,0.0000,-1039.9,-1498.5,-735.56,-1149.1
1861.000000000,73.588,1710.2,1748.3,1762.7,259.83,3970.3,966.86,2.6041,6274.4,2754.4,3375.9,2105.1,0.0000,-5754.4,-6487.2,-992.04,-1755.8,-1425.1,-14775.,-88.527,-18573.,-5945.6,-3819.3,-2082.5,55.500,1977.2,1802.8,1799.6,285.57,4122.9,1686.6,0.0000,7306.6,4449.7,4252.8,3658.0,0.0000,-288.07,-87.495,-88.085,-37.000,-98.123,-587.69,0.0000,-1039.9,-1498.4,-735.54,-1149.0
1862.000000000,73.459,1706.3,1744.0,1751.6,259.10,3944.6,966.86,2.6045,6259.0,2754.4,3376.0,2105.2,0.0000,-5750.6,-6485.4,-990.96,-1755.2,-1424.1,-14774.,-88.502,-18572.,-5945.2,-3819.1,-2082.1,55.361,1972.2,1798.3,1787.5,284.72,4092.8,1686.6,0.0000,7288.3,4449.7,4252.8,3658.0,0.0000,-287.26,-87.248,-87.604,-36.907,-97.377,-587.69,0.0000,-1039.9,-1498.4,-735.52,-1148.9
1863.000000000,73.322,1702.6,1739.9,1740.3,258.38,3918.8,966.86,2.6049,6243.5,2754.5,3376.0,2105.3,0.0000,-5746.7,-6483.7,-989.82,-1754.5,-1423.0,-14774.,-88.476,-18572.,-5944.9,-3818.9,-2081.7,55.236,1967.8,1794.3,1775.8,283.95,4063.9,1686.6,0.0000,7270.8,4449.7,4252.8,3658.0,0.0000,-286.53,-87.025,-87.146,-36.824,-96.656,-587.69,0.0000,-1039.9,-1498.3,-735.50,-1148.8
1864.000000000,73.197,1699.2,1736.0,1729.2,257.68,3893.2,966.86,2.6053,6227.9,2754.6,3376.0,2105.5,0.0000,-5742.8,-6481.9,-988.64,-1753.8,-1421.7,-14773.,-88.451,-18571.,-5944.5,-3818.7,-2081.3,55.133,1964.1,1790.9,1764.6,283.28,4036.1,1686.6,0.0000,7253.9,4449.7,4252.8,3658.0,0.0000,-285.91,-86.835,-86.717,-36.755,-95.958,-587.69,0.0000,-1039.9,-1498.3,-735.48,-1148.7
1865.000000000,73.076,1695.7,1732.5,1718.4,257.02,3876.8,966.86,2.6057,6212.2,2754.6,3375.9,2105.6,0.0000,-5738.9,-6480.1,-987.41,-1753.1,-1420.4,-14772.,-88.425,-18570.,-5944.2,-3818.4,-2080.9,55.029,1960.4,1787.5,1753.7,282.62,4008.9,1686.6,0.0000,7237.3,4449.7,4252.8,3658.0,0.0000,-285.28,-86.645,-86.294,-36.686,-95.272,-587.69,0.0000,-1039.9,-1498.2,-735.46,-1148.6
1866.000000000,72.935,1692.1,1729.0,1707.7,256.41,3852.5,966.86,2.6061,6196.4,2754.7,3375.8,2105.7,0.0000,-5735.0,-6478.4,-986.14,-1752.5,-1418.9,-14771.,-88.400,-18569.,-5943.8,-3818.2,-2080.5,54.913,1956.3,1783.8,1742.5,281.90,3981.1,1686.6,0.0000,7220.5,4449.7,4252.8,3658.0,0.0000,-284.60,-86.436,-85.857,-36.609,-94.572,-587.69,0.0000,-1039.9,-1498.2,-735.43,-1148.5
1867.000000000,72.817,1688.7,1725.6,1697.1,255.78,3827.3,966.86,2.6065,6180.6,2754.7,3375.9,2105.8,0.0000,-5731.1,-6476.6,-984.83,-1751.8,-1417.4,-14771.,-88.374,-18569.,-5943.5,-3818.0,-2080.1,54.782,1951.6,1779.5,1731.0,281.09,3952.7,1686.6,0.0000,7203.2,4449.7,4252.8,3658.0,0.0000,-283.83,-86.202,-85.400,-36.521,-93.853,-587.69,0.0000,-1039.9,-1498.1,-735.41,-1148.4
1868.000000000,72.698,1685.1,1722.0,1686.6,255.09,3801.9,966.86,2.6069,6164.7,2754.8,3376.0,2105.9,0.0000,-5727.1,-6474.9,-983.48,-1751.1,-1415.7,-14770.,-88.349,-18568.,-5943.2,-3817.8,-2079.7,54.666,1947.4,1775.7,1719.9,280.37,3925.2,1686.6,0.0000,7186.6,4449.7,4252.8,3658.0,0.0000,-283.14,-85.992,-84.965,-36.444,-93.155,-587.69,0.0000,-1039.9,-1498.0,-735.39,-1148.3
1869.000000000,72.581,1681.6,1718.4,1676.2,254.42,3776.6,966.86,2.6073,6149.0,2754.8,3376.0,2106.0,0.0000,-5723.2,-6473.1,-982.09,-1750.4,-1413.9,-14769.,-88.323,-18567.,-5942.8,-3817.6,-2079.3,54.572,1944.1,1772.7,1709.6,279.76,3899.3,1686.6,0.0000,7170.8,4449.7,4252.8,3658.0,0.0000,-282.56,-85.817,-84.565,-36.381,-92.492,-587.69,0.0000,-1039.9,-1498.0,-735.37,-1148.2
1870.000000000,72.472,1678.6,1715.1,1665.9,253.84,3751.8,966.86,2.6077,6133.6,2754.9,3376.1,2106.1,0.0000,-5719.3,-6471.3,-980.68,-1749.8,-1412.0,-14768.,-88.298,-18566.,-5942.5,-3817.3,-2078.9,54.509,1941.9,1770.7,1700.5,279.32,3876.6,1686.6,0.0000,7157.0,4449.7,4252.8,3658.0,0.0000,-282.15,-85.693,-84.225,-36.340,-91.905,-587.69,0.0000,-1039.9,-1497.9,-735.35,-1148.2
1871.000000000,72.376,1675.9,1712.3,1656.0,253.31,3727.6,966.86,2.6081,6118.6,2754.9,3376.1,2106.2,0.0000,-5715.4,-6469.6,-979.24,-1749.1,-1410.1,-14768.,-88.273,-18565.,-5942.1,-3817.1,-2078.5,54.397,1937.9,1767.0,1690.0,278.62,3850.4,1686.6,0.0000,7141.1,4449.7,4252.8,3658.0,0.0000,-281.48,-85.489,-83.809,-36.264,-91.233,-587.69,0.0000,-1039.9,-1497.9,-735.32,-1148.1
1872.000000000,72.277,1672.7,1709.2,1646.3,252.70,3703.6,966.86,2.6085,6103.7,2755.0,3376.1,2106.3,0.0000,-5711.5,-6467.9,-977.76,-1748.4,-1408.1,-14767.,-88.247,-18564.,-5941.8,-3816.9,-2078.1,54.245,1932.5,1762.1,1678.4,277.73,3821.9,1686.6,0.0000,7123.8,4449.7,4252.8,3658.0,0.0000,-280.61,-85.225,-83.337,-36.164,-90.503,-587.69,0.0000,-1039.9,-1497.8,-735.30,-1148.0
1873.000000000,72.200,1668.6,1705.4,1636.4,252.02,3679.1,966.86,2.6088,6088.7,2755.0,3376.0,2106.4,0.0000,-5707.6,-6466.2,-976.25,-1747.7,-1406.0,-14766.,-88.222,-18563.,-5941.5,-3816.7,-2077.7,54.092,1927.0,1757.1,1666.7,276.83,3793.5,1686.6,0.0000,7106.6,4449.7,4252.8,3658.0,0.0000,-279.73,-84.957,-82.865,-36.061,-89.773,-587.69,0.0000,-1040.0,-1497.8,-735.28,-1147.9
1874.000000000,72.107,1664.6,1701.3,1626.3,251.31,3654.1,966.86,2.6093,6073.5,2755.3,3376.0,2106.5,0.0000,-5703.6,-6464.4,-974.71,-1747.1,-1403.7,-14765.,-88.197,-18562.,-5941.1,-3816.4,-2077.3,53.948,1921.9,1752.4,1655.4,275.97,3765.6,1686.6,0.0000,7089.6,4449.7,4252.8,3658.0,0.0000,-278.89,-84.703,-82.406,-35.965,-89.055,-587.69,0.0000,-1040.0,-1497.7,-735.26,-1147.8
1875.000000000,72.078,1660.5,1697.1,1616.0,250.55,3629.0,966.83,2.6096,6058.4,2755.4,3376.1,2106.6,0.0000,-5699.5,-6462.6,-973.13,-1746.4,-1401.4,-14764.,-88.171,-18561.,-5940.8,-3816.2,-2076.9,53.797,1916.5,1747.5,1643.9,275.08,3737.6,1686.6,0.0000,7072.6,4449.7,4252.8,3658.0,0.0000,-278.03,-84.439,-81.940,-35.865,-88.332,-587.69,0.0000,-1040.0,-1497.7,-735.24,-1147.7
1876.000000000,72.003,1656.5,1693.1,1605.6,249.80,3604.1,966.82,2.6100,6043.4,2755.5,3376.0,2106.8,0.0000,-5695.5,-6460.7,-971.52,-1745.7,-1399.0,-14763.,-88.146,-18559.,-5940.5,-3816.0,-2076.5,53.712,1913.5,1744.8,1634.2,274.53,3713.3,1686.6,0.0000,7057.9,4449.7,4252.8,3658.0,0.0000,-277.50,-84.279,-81.566,-35.808,-87.698,-587.69,0.0000,-1040.0,-1497.6,-735.21,-1147.6
1877.000000000,71.876,1654.2,1690.3,1595.5,249.34,3580.3,966.82,2.6104,6028.8,2755.5,3375.9,2106.8,0.0000,-5691.5,-6458.9,-969.90,-1745.0,-1396.6,-14762.,-88.121,-18558.,-5940.1,-3815.8,-2076.1,54.138,1919.8,1750.5,1629.3,275.24,3698.5,1686.6,0.58015E-02,7048.8,4449.7,4252.9,3658.1,0.0000,-278.31,-84.528,-81.480,-35.924,-87.286,-587.69,-0.26489E-03,-1040.0,-1497.6,-735.19,-1147.5
1878.000000000,71.888,1659.2,1694.3,1587.1,250.09,3560.5,966.82,2.6108,6014.9,2755.6,3375.9,2106.9,0.0000,-5688.0,-6457.5,-968.40,-1744.3,-1394.2,-14761.,-88.099,-18557.,-5939.8,-3815.5,-2075.8,63.995,1971.5,1800.0,1655.6,281.96,3750.2,1686.6,2.1173,7079.8,4450.7,4255.2,3659.8,0.0000,-284.92,-86.698,-82.945,-36.789,-88.428,-587.69,-0.96675E-01,-1040.0,-1497.5,-735.18,-1147.4
1879.000000000,72.360,1675.9,1708.7,1583.5,252.79,3548.5,966.82,2.6112,6002.9,2755.6,3375.9,2107.1,0.0000,-5685.7,-6456.9,-967.02,-1743.9,-1391.9,-14760.,-88.076,-18556.,-5939.5,-3815.3,-2075.4,55.819,1988.5,1813.2,1651.3,284.96,3735.2,1686.6,0.0000,7071.2,4451.4,4254.6,3658.5,0.0000,-288.14,-87.526,-83.176,-37.215,-88.027,-587.69,0.0000,-1040.0,-1497.5,-735.16,-1147.3
1880.000000000,72.969,1691.4,1723.7,1583.9,254.66,3538.8,966.82,2.6116,5992.2,2755.7,3375.9,2107.1,0.0000,-5684.3,-6456.9,-965.68,-1743.5,-1390.0,-14760.,-88.053,-18554.,-5939.1,-3815.1,-2075.0,55.937,1992.7,1817.0,1642.6,285.31,3711.2,1686.6,0.0000,7056.7,4451.3,4254.5,3658.5,0.0000,-288.69,-87.702,-82.944,-37.294,-87.406,-587.69,0.0000,-1040.0,-1497.4,-735.13,-1147.2
1881.000000000,73.303,1699.8,1732.3,1582.5,255.99,3525.0,966.82,2.6120,5980.9,2755.7,3376.0,2107.2,0.0000,-5683.1,-6457.0,-964.39,-1743.2,-1387.9,-14759.,-88.029,-18553.,-5938.8,-3814.8,-2074.6,55.952,1993.3,1817.5,1633.1,285.13,3685.8,1686.6,0.0000,7041.0,4450.6,4253.9,3658.3,0.0000,-288.71,-87.718,-82.631,-37.304,-86.761,-587.69,0.0000,-1040.0,-1497.4,-735.11,-1147.1
1882.000000000,73.756,1703.6,1736.0,1579.7,257.09,3507.9,966.82,2.6111,5968.9,2755.8,3375.9,2107.3,0.0000,-5682.0,-6457.0,-963.10,-1742.8,-1385.7,-14758.,-88.005,-18552.,-5938.5,-3814.6,-2074.2,55.879,1990.7,1815.1,1622.5,284.47,3658.9,1686.6,0.0000,7024.5,4450.2,4253.4,3658.2,0.0000,-288.27,-87.594,-82.239,-37.254,-86.075,-587.69,0.0000,-1040.0,-1497.3,-735.08,-1147.0
1883.000000000,73.970,1704.2,1737.5,1573.8,257.17,3488.7,966.82,2.6076,5958.5,2755.9,3375.9,2107.4,0.0000,-5680.8,-6456.9,-961.86,-1742.4,-1383.4,-14757.,-87.980,-18550.,-5938.1,-3814.4,-2073.8,55.783,1987.2,1812.0,1612.0,283.75,3632.4,1686.6,0.0000,7008.3,4449.9,4253.1,3658.1,0.0000,-287.72,-87.435,-81.836,-37.189,-85.396,-587.69,0.0000,-1040.0,-1497.3,-735.06,-1146.9
1884.000000000,73.953,1703.4,1737.0,1566.0,256.80,3468.9,966.82,2.6080,5949.8,2755.9,3375.9,2107.5,0.0000,-5679.5,-6456.7,-960.51,-1741.9,-1380.9,-14756.,-87.955,-18549.,-5937.8,-3814.1,-2073.4,55.671,1983.3,1808.4,1601.5,283.00,3606.3,1686.6,0.0000,6992.4,4449.8,4252.9,3658.0,0.0000,-287.08,-87.250,-81.425,-37.114,-84.723,-587.69,0.0000,-1040.0,-1497.2,-735.04,-1146.8
1885.000000000,73.886,1701.6,1735.5,1557.1,256.27,3453.1,966.78,2.6084,5944.2,2756.0,3375.8,2107.5,0.0000,-5677.9,-6456.3,-959.06,-1741.4,-1378.3,-14755.,-87.930,-18548.,-5937.5,-3813.9,-2073.0,55.525,1978.1,1803.7,1590.6,282.12,3579.4,1686.6,0.0000,6976.1,4449.7,4252.8,3658.0,0.0000,-286.27,-87.011,-80.980,-37.017,-84.027,-587.69,0.0000,-1040.0,-1497.2,-735.01,-1146.7
1886.000000000,73.773,1698.9,1734.2,1547.8,255.64,3438.1,966.74,2.6132,5936.1,2756.2,3375.8,2107.6,0.0000,-5676.2,-6455.7,-957.55,-1740.9,-1375.6,-14754.,-87.905,-18546.,-5937.1,-3813.6,-2072.6,55.449,1975.3,1801.2,1581.4,281.60,3556.4,1686.6,0.0000,6962.1,4449.7,4252.8,3658.0,0.0000,-285.82,-86.880,-80.629,-36.966,-83.422,-587.69,0.0000,-1040.0,-1497.1,-734.99,-1146.6
1887.000000000,73.668,1697.3,1733.0,1538.6,255.07,3419.3,966.74,2.6138,5925.2,2756.3,3375.9,2107.7,0.0000,-5674.4,-6455.2,-955.98,-1740.4,-1372.9,-14753.,-87.880,-18545.,-5936.8,-3813.4,-2072.2,55.317,1970.6,1796.9,1571.2,280.82,3531.4,1686.6,0.0000,6947.0,4449.7,4252.8,3658.0,0.0000,-285.08,-86.661,-80.215,-36.878,-82.767,-587.69,0.0000,-1040.0,-1497.1,-734.97,-1146.5
1888.000000000,73.558,1695.3,1730.9,1530.5,254.42,3397.9,966.74,2.6141,5912.3,2756.4,3375.9,2107.8,0.0000,-5672.4,-6454.5,-954.37,-1739.9,-1370.0,-14752.,-87.855,-18543.,-5936.5,-3813.1,-2071.8,55.175,1965.6,1792.3,1560.9,279.99,3506.3,1686.6,0.0000,6931.7,4449.7,4252.8,3658.0,0.0000,-284.29,-86.425,-79.793,-36.784,-82.109,-587.69,0.0000,-1040.0,-1497.0,-734.95,-1146.4
1889.000000000,73.416,1691.9,1727.2,1521.9,253.72,3375.1,966.74,2.6145,5898.4,2756.4,3375.8,2107.9,0.0000,-5670.3,-6453.7,-952.73,-1739.4,-1367.2,-14751.,-87.830,-18542.,-5936.2,-3812.9,-2071.4,55.017,1959.9,1787.1,1550.4,279.08,3480.7,1686.6,0.0000,6916.2,4449.7,4252.8,3658.0,0.0000,-283.41,-86.162,-79.354,-36.678,-81.437,-587.69,0.0000,-1040.0,-1497.0,-734.93,-1146.3
1890.000000000,73.289,1688.4,1722.9,1512.6,252.98,3352.6,966.70,2.6166,5884.2,2756.5,3375.8,2108.0,0.0000,-5667.9,-6452.8,-951.04,-1738.8,-1364.2,-14749.,-87.805,-18541.,-5935.8,-3812.7,-2071.0,54.836,1953.5,1781.3,1539.4,278.06,3454.3,1686.6,0.0000,6900.2,4449.7,4252.8,3658.0,0.0000,-282.42,-85.862,-78.890,-36.557,-80.746,-587.69,0.0000,-1040.0,-1496.9,-734.90,-1146.2
1891.000000000,73.130,1684.9,1719.0,1502.9,252.17,3330.5,966.70,2.6431,5870.6,2756.5,3375.7,2108.1,0.0000,-5665.4,-6451.9,-949.33,-1738.3,-1361.3,-14748.,-87.780,-18539.,-5935.5,-3812.4,-2070.6,54.679,1947.9,1776.2,1529.1,277.17,3429.3,1686.6,0.0000,6885.0,4449.7,4252.8,3658.0,0.0000,-281.54,-85.600,-78.460,-36.453,-80.090,-587.69,0.0000,-1040.0,-1496.9,-734.88,-1146.1
1892.000000000,72.970,1681.0,1715.3,1493.2,251.41,3308.9,966.71,2.6434,5857.1,2756.6,3375.8,2108.2,0.0000,-5662.6,-6450.8,-947.59,-1737.7,-1358.2,-14747.,-87.755,-18538.,-5935.2,-3812.2,-2070.2,54.532,1942.7,1771.4,1519.2,276.32,3405.1,1686.6,0.0000,6870.3,4449.7,4252.8,3658.0,0.0000,-280.72,-85.352,-78.046,-36.355,-79.450,-587.69,0.0000,-1040.0,-1496.8,-734.86,-1146.0
1893.000000000,72.889,1677.1,1711.2,1483.9,250.63,3286.8,966.71,2.6438,5843.1,2756.6,3375.8,2108.4,0.0000,-5659.8,-6449.7,-945.81,-1737.1,-1355.2,-14746.,-87.730,-18536.,-5934.8,-3811.9,-2069.8,54.390,1937.6,1766.8,1509.4,275.50,3381.4,1686.6,0.0000,6855.9,4449.7,4252.8,3658.0,0.0000,-279.92,-85.111,-77.641,-36.260,-78.820,-587.69,0.0000,-1040.0,-1496.8,-734.84,-1145.9
1894.000000000,72.758,1673.4,1707.4,1474.5,249.86,3264.6,966.71,2.6441,5829.4,2756.7,3375.9,2108.4,0.0000,-5656.9,-6448.6,-944.01,-1736.5,-1352.0,-14745.,-87.705,-18534.,-5934.5,-3811.7,-2069.4,54.236,1932.1,1761.8,1499.5,274.63,3357.3,1686.6,0.0000,6841.3,4449.7,4252.8,3658.0,0.0000,-279.06,-84.852,-77.224,-36.158,-78.182,-587.69,0.0000,-1040.0,-1496.7,-734.81,-1145.8
1895.000000000,72.606,1669.3,1703.9,1465.1,249.08,3242.3,966.71,2.6445,5816.0,2756.7,3376.0,2108.5,0.0000,-5653.9,-6447.4,-942.17,-1735.9,-1348.8,-14744.,-87.680,-18533.,-5934.2,-3811.4,-2069.0,54.063,1926.0,1756.2,1489.2,273.66,3332.5,1686.6,0.0000,6826.3,4449.7,4252.8,3658.0,0.0000,-278.10,-84.561,-76.785,-36.042,-77.526,-587.69,0.0000,-1040.0,-1496.7,-734.79,-1145.8
1896.000000000,72.446,1664.9,1699.5,1455.6,248.20,3220.4,966.71,2.6449,5802.3,2756.8,3376.0,2108.6,0.0000,-5650.9,-6446.1,-940.31,-1735.3,-1345.6,-14743.,-87.655,-18531.,-5933.8,-3811.2,-2068.6,53.862,1918.8,1749.6,1478.3,272.54,3306.5,1686.6,0.0000,6810.5,4449.7,4252.8,3658.0,0.0000,-276.99,-84.225,-76.312,-35.908,-76.841,-587.69,0.0000,-1040.0,-1496.6,-734.77,-1145.7
1897.000000000,72.324,1660.2,1694.5,1446.1,247.34,3198.0,966.71,2.6452,5788.5,2756.9,3376.0,2108.7,0.0000,-5647.7,-6444.7,-938.42,-1734.7,-1342.4,-14742.,-87.630,-18530.,-5933.5,-3810.9,-2068.2,53.716,1913.6,1744.9,1468.8,271.71,3283.3,1686.6,0.0000,6796.4,4449.7,4252.8,3658.0,0.0000,-276.16,-83.975,-75.911,-35.810,-76.224,-587.69,0.0000,-1040.0,-1496.6,-734.75,-1145.6
1898.000000000,72.088,1655.8,1689.5,1436.5,246.56,3175.9,966.71,2.6303,5774.7,2757.2,3376.1,2108.8,0.0000,-5644.4,-6443.3,-936.51,-1734.1,-1339.0,-14741.,-87.605,-18528.,-5933.2,-3810.7,-2067.8,53.570,1908.4,1740.1,1459.3,270.88,3260.4,1686.6,0.0000,6782.5,4449.7,4252.8,3658.0,0.0000,-275.34,-83.724,-75.514,-35.713,-75.612,-587.69,0.0000,-1040.0,-1496.5,-734.72,-1145.5
1899.000000000,71.919,1651.2,1684.9,1427.1,245.78,3154.2,966.71,2.5789,5761.6,2757.3,3376.2,2108.8,0.0000,-5641.0,-6441.8,-934.58,-1733.4,-1335.7,-14740.,-87.580,-18526.,-5932.9,-3810.4,-2067.4,53.419,1903.0,1735.2,1449.8,270.02,3237.4,1686.6,0.0000,6768.5,4449.7,4252.8,3658.0,0.0000,-274.49,-83.467,-75.112,-35.613,-74.997,-587.69,0.0000,-1040.0,-1496.5,-734.70,-1145.4
1900.000000000,71.807,1646.8,1680.6,1417.8,245.00,3132.7,966.70,2.5792,5748.9,2757.3,3376.2,2108.8,0.0000,-5637.6,-6440.3,-932.63,-1732.8,-1332.2,-14738.,-87.555,-18525.,-5932.5,-3810.1,-2067.0,53.268,1897.6,1730.3,1440.3,269.17,3214.5,1686.6,0.0000,6754.7,4449.7,4252.8,3658.0,0.0000,-273.64,-83.208,-74.712,-35.512,-74.386,-587.69,0.0000,-1040.0,-1496.4,-734.68,-1145.3
1901.000000000,71.655,1642.4,1676.0,1408.9,244.23,3111.4,966.68,2.5796,5735.9,2757.4,3376.2,2108.9,0.0000,-5634.1,-6438.8,-930.65,-1732.1,-1328.8,-14737.,-87.530,-18523.,-5932.2,-3809.9,-2066.7,53.098,1891.6,1724.8,1430.5,268.22,3191.0,1686.6,0.0000,6740.4,4449.7,4252.8,3658.0,0.0000,-272.68,-82.919,-74.291,-35.399,-73.758,-587.69,0.0000,-1040.0,-1496.3,-734.66,-1145.2
1902.000000000,71.498,1638.0,1671.2,1399.8,243.41,3090.4,966.64,2.5799,5722.8,2757.4,3376.3,2109.0,0.0000,-5630.5,-6437.2,-928.66,-1731.5,-1325.3,-14736.,-87.505,-18521.,-5931.9,-3809.6,-2066.3,52.916,1885.1,1718.9,1420.5,267.21,3166.9,1686.6,0.0000,6725.8,4449.7,4252.8,3658.0,0.0000,-271.67,-82.609,-73.855,-35.277,-73.118,-587.69,0.0000,-1039.9,-1496.3,-734.63,-1145.1
1903.000000000,71.330,1633.1,1666.1,1390.9,242.56,3069.1,966.64,2.5803,5709.3,2757.5,3376.3,2109.1,0.0000,-5626.7,-6435.5,-926.64,-1730.8,-1321.7,-14735.,-87.480,-18520.,-5931.6,-3809.4,-2065.9,52.726,1878.3,1712.7,1410.3,266.17,3142.7,1686.6,0.0000,6711.1,4449.7,4252.8,3658.0,0.0000,-270.61,-82.289,-73.413,-35.151,-72.474,-587.69,0.0000,-1039.9,-1496.2,-734.61,-1145.0
1904.000000000,70.885,1627.8,1660.9,1381.8,241.69,3047.1,966.64,2.5806,5695.8,2757.5,3376.3,2109.1,0.0000,-5622.9,-6433.7,-924.60,-1730.1,-1318.2,-14734.,-87.455,-18518.,-5931.2,-3809.1,-2065.5,52.538,1871.7,1706.6,1400.3,265.13,3118.6,1686.6,0.0000,6696.5,4449.7,4252.8,3658.0,0.0000,-269.57,-81.970,-72.975,-35.026,-71.835,-587.69,0.0000,-1039.9,-1496.2,-734.59,-1144.9
1905.000000000,70.703,1622.3,1656.4,1372.5,240.81,3025.5,966.64,2.5810,5682.4,2757.3,3376.3,2109.2,0.0000,-5619.1,-6432.0,-922.54,-1729.4,-1314.5,-14732.,-87.431,-18516.,-5930.9,-3808.8,-2065.1,52.381,1866.0,1701.5,1390.9,264.25,3096.2,1686.6,0.0000,6682.9,4449.7,4252.8,3658.0,0.0000,-268.67,-81.698,-72.576,-34.920,-71.234,-587.69,0.0000,-1039.9,-1496.1,-734.57,-1144.8
1906.000000000,70.527,1617.6,1652.2,1363.3,239.98,3004.3,966.64,2.5813,5669.2,2757.4,3376.3,2109.3,0.0000,-5615.2,-6430.1,-920.47,-1728.7,-1310.8,-14731.,-87.406,-18514.,-5930.6,-3808.6,-2064.7,52.230,1860.7,1696.6,1381.8,263.40,3074.3,1686.6,0.0000,6669.6,4449.7,4252.8,3658.0,0.0000,-267.82,-81.436,-72.188,-34.820,-70.643,-587.69,0.0000,-1039.9,-1496.1,-734.54,-1144.7
1907.000000000,70.360,1613.0,1647.5,1354.1,239.17,2983.6,966.64,2.5816,5656.1,2757.4,3376.4,2109.4,0.0000,-5611.3,-6428.3,-918.37,-1728.0,-1307.1,-14730.,-87.381,-18513.,-5930.3,-3808.3,-2064.3,52.065,1854.8,1691.3,1372.5,262.49,3051.8,1686.6,0.0000,6656.0,4449.7,4252.8,3658.0,0.0000,-266.89,-81.153,-71.785,-34.710,-70.042,-587.69,0.0000,-1039.9,-1496.0,-734.52,-1144.6
1908.000000000,70.192,1608.2,1642.6,1345.3,238.35,2963.0,966.64,2.5820,5643.1,2757.5,3376.4,2109.5,0.0000,-5607.3,-6426.4,-916.26,-1727.3,-1303.3,-14729.,-87.356,-18511.,-5929.9,-3808.0,-2063.9,51.887,1848.5,1685.5,1362.9,261.50,3028.9,1686.6,0.0000,6642.1,4449.7,4252.8,3658.0,0.0000,-265.89,-80.848,-71.367,-34.591,-69.428,-587.69,0.0000,-1039.9,-1496.0,-734.50,-1144.5
1909.000000000,70.023,1603.1,1637.8,1336.6,237.53,2942.2,966.64,2.5823,5630.2,2757.5,3376.4,2109.5,0.0000,-5603.2,-6424.5,-914.14,-1726.6,-1299.5,-14728.,-87.331,-18509.,-5929.6,-3807.8,-2063.5,51.702,1841.9,1679.5,1353.2,260.49,3005.8,1686.6,0.0000,6628.1,4449.7,4252.8,3658.0,0.0000,-264.86,-80.533,-70.942,-34.468,-68.812,-587.69,0.0000,-1039.9,-1495.9,-734.47,-1144.4
1910.000000000,69.850,1597.9,1633.0,1327.8,236.68,2921.2,966.64,2.5827,5617.4,2757.6,3376.4,2109.6,0.0000,-5599.2,-6422.6,-911.99,-1725.9,-1295.6,-14726.,-87.307,-18507.,-5929.3,-3807.5,-2063.1,51.507,1834.9,1673.1,1343.3,259.42,2982.4,1686.6,0.0000,6613.9,4449.7,4252.8,3658.0,0.0000,-263.77,-80.201,-70.507,-34.338,-68.187,-587.69,0.0000,-1039.9,-1495.9,-734.45,-1144.3
1911.000000000,69.669,1592.4,1627.6,1318.8,235.78,2900.1,966.64,2.5830,5604.3,2757.6,3376.5,2109.6,0.0000,-5595.0,-6420.6,-909.83,-1725.1,-1291.7,-14725.,-87.282,-18506.,-5929.0,-3807.2,-2062.7,51.310,1827.9,1666.7,1333.5,258.35,2959.0,1686.6,0.0000,6599.7,4449.7,4252.8,3658.0,0.0000,-262.66,-79.865,-70.071,-34.206,-67.565,-587.69,0.0000,-1039.9,-1495.8,-734.43,-1144.2
1912.000000000,69.274,1586.9,1622.0,1309.7,234.87,2879.3,966.64,2.5834,5591.4,2757.7,3376.5,2109.7,0.0000,-5590.7,-6418.5,-907.65,-1724.4,-1287.7,-14724.,-87.257,-18504.,-5928.6,-3807.0,-2062.3,51.125,1821.3,1660.7,1324.0,257.34,2936.4,1686.6,0.0000,6586.0,4449.7,4252.8,3658.0,0.0000,-261.63,-79.549,-69.653,-34.084,-66.959,-587.69,0.0000,-1039.9,-1495.8,-734.41,-1144.1
1913.000000000,69.010,1581.8,1616.7,1300.7,234.02,2858.4,966.64,2.5698,5578.6,2757.7,3376.5,2109.8,0.0000,-5586.4,-6416.4,-905.46,-1723.7,-1283.7,-14722.,-87.232,-18502.,-5928.3,-3806.7,-2061.9,51.044,1818.4,1658.1,1316.0,256.83,2916.7,1686.6,0.0000,6574.0,4449.7,4252.8,3658.0,0.0000,-261.13,-79.394,-69.340,-34.029,-66.423,-587.69,0.0000,-1039.9,-1495.7,-734.38,-1144.0
1914.000000000,68.837,1577.7,1612.1,1291.7,233.25,2837.9,966.64,2.5507,5565.9,2757.8,3376.5,2109.8,0.0000,-5582.0,-6414.4,-903.26,-1722.9,-1279.7,-14721.,-87.208,-18500.,-5928.0,-3806.4,-2061.5,50.894,1813.1,1653.2,1307.4,255.99,2896.0,1686.6,0.0000,6561.5,4449.7,4252.8,3658.0,0.0000,-260.27,-79.132,-68.968,-33.929,-65.862,-587.69,0.0000,-1039.9,-1495.7,-734.36,-1143.9
1915.000000000,68.648,1573.4,1607.7,1283.1,232.44,2817.8,966.64,2.5510,5553.6,2757.8,3376.5,2109.8,0.0000,-5577.7,-6412.4,-901.05,-1722.2,-1275.6,-14720.,-87.183,-18498.,-5927.7,-3806.1,-2061.1,50.737,1807.5,1648.1,1298.7,255.13,2875.0,1686.6,0.0000,6548.8,4449.7,4252.8,3658.0,0.0000,-259.37,-78.860,-68.590,-33.825,-65.297,-587.69,0.0000,-1039.9,-1495.6,-734.34,-1143.8
1916.000000000,68.483,1568.9,1603.2,1274.7,231.70,2797.9,966.64,2.5514,5541.5,2757.9,3376.5,2109.9,0.0000,-5573.3,-6410.3,-898.83,-1721.4,-1271.5,-14719.,-87.159,-18496.,-5927.3,-3805.9,-2060.7,50.576,1801.7,1642.9,1289.9,254.24,2854.0,1686.6,0.0000,6536.0,4449.7,4252.8,3658.0,0.0000,-258.46,-78.580,-68.208,-33.717,-64.731,-587.69,0.0000,-1039.9,-1495.6,-734.31,-1143.7
1917.000000000,68.209,1564.2,1598.2,1266.4,230.98,2778.1,966.62,2.5517,5529.1,2757.9,3376.4,2110.0,0.0000,-5568.8,-6408.3,-896.60,-1720.7,-1267.4,-14717.,-87.134,-18494.,-5927.0,-3805.6,-2060.3,50.399,1795.4,1637.1,1280.8,253.27,2832.5,1686.6,0.0000,6522.9,4449.7,4252.8,3658.0,0.0000,-257.46,-78.276,-67.809,-33.599,-64.152,-587.69,0.0000,-1039.8,-1495.5,-734.29,-1143.6
1918.000000000,67.995,1559.2,1593.0,1258.0,230.17,2758.2,966.62,2.5520,5516.6,2758.0,3376.4,2110.2,0.0000,-5564.3,-6406.2,-894.36,-1719.9,-1263.3,-14716.,-87.109,-18492.,-5926.7,-3805.3,-2059.9,50.226,1789.3,1631.5,1271.9,252.32,2811.2,1686.6,0.0000,6510.0,4449.7,4252.8,3658.0,0.0000,-256.48,-77.977,-67.415,-33.484,-63.579,-587.69,0.0000,-1039.8,-1495.5,-734.27,-1143.5
1919.000000000,67.825,1554.1,1587.7,1249.5,229.36,2738.4,966.62,2.5523,5504.2,2758.0,3376.5,2110.3,0.0000,-5559.8,-6404.1,-892.11,-1719.1,-1259.1,-14715.,-87.085,-18490.,-5926.4,-3805.0,-2059.6,50.050,1783.0,1625.8,1262.9,251.36,2789.9,1686.6,0.0000,6497.1,4449.7,4252.8,3658.0,0.0000,-255.49,-77.675,-67.020,-33.366,-63.008,-587.69,0.0000,-1039.8,-1495.4,-734.25,-1143.4
1920.000000000,67.655,1549.0,1582.3,1241.4,228.56,2718.5,966.62,2.5527,5491.9,2758.1,3376.4,2110.3,0.0000,-5555.1,-6401.9,-889.85,-1718.4,-1254.9,-14713.,-87.060,-18488.,-5926.1,-3804.7,-2059.2,49.880,1777.0,1620.3,1254.1,250.43,2769.0,1686.6,0.0000,6484.5,4449.7,4252.8,3658.0,0.0000,-254.53,-77.382,-66.635,-33.254,-62.446,-587.69,0.0000,-1039.8,-1495.4,-734.22,-1143.3
1921.000000000,67.481,1543.9,1576.9,1233.1,227.74,2698.7,966.62,2.5530,5479.8,2758.1,3376.4,2110.4,0.0000,-5550.5,-6399.8,-887.58,-1717.6,-1250.7,-14712.,-87.035,-18486.,-5925.7,-3804.5,-2058.8,49.735,1771.8,1615.6,1245.9,249.62,2749.3,1686.6,0.0000,6472.5,4449.7,4252.8,3658.0,0.0000,-253.69,-77.127,-66.280,-33.156,-61.912,-587.69,0.0000,-1039.8,-1495.3,-734.20,-1143.2
1922.000000000,67.317,1539.1,1572.0,1224.7,226.95,2679.5,966.62,2.5533,5467.8,2758.2,3376.5,2110.5,0.0000,-5545.7,-6397.6,-885.30,-1716.8,-1246.4,-14710.,-87.011,-18484.,-5925.4,-3804.2,-2058.4,49.571,1766.0,1610.3,1237.4,248.73,2729.0,1686.6,0.0000,6460.2,4449.7,4252.8,3658.0,0.0000,-252.76,-76.843,-65.906,-33.048,-61.365,-587.69,0.0000,-1039.8,-1495.3,-734.18,-1143.2
1923.000000000,67.155,1534.4,1567.1,1216.4,226.15,2660.6,966.62,2.5536,5456.0,2758.2,3376.5,2110.6,0.0000,-5541.0,-6395.4,-883.02,-1716.0,-1242.1,-14709.,-86.986,-18482.,-5925.1,-3803.9,-2058.0,49.414,1760.3,1605.1,1229.0,247.86,2709.0,1686.6,0.0000,6448.1,4449.7,4252.8,3658.0,0.0000,-251.86,-76.569,-65.540,-32.942,-60.825,-587.69,0.0000,-1039.8,-1495.2,-734.15,-1143.1
1924.000000000,66.990,1529.7,1562.3,1208.5,225.41,2641.8,966.62,2.5540,5444.4,2758.3,3376.6,2110.7,0.0000,-5536.3,-6393.3,-880.73,-1715.2,-1237.8,-14708.,-86.962,-18480.,-5924.8,-3803.6,-2057.6,49.305,1756.5,1601.6,1221.7,247.23,2691.3,1686.6,0.0000,6437.3,4449.7,4252.8,3658.0,0.0000,-251.21,-76.370,-65.235,-32.870,-60.338,-587.69,0.0000,-1039.8,-1495.2,-734.13,-1143.0
1925.000000000,66.847,1525.5,1557.8,1200.7,224.75,2623.1,966.62,2.5543,5432.7,2758.3,3376.6,2110.8,0.0000,-5531.5,-6391.1,-878.44,-1714.4,-1233.5,-14706.,-86.937,-18478.,-5924.5,-3803.3,-2057.2,49.160,1751.3,1596.9,1213.7,246.43,2672.2,1686.6,0.0000,6425.7,4449.7,4252.8,3658.0,0.0000,-250.38,-76.117,-64.889,-32.774,-59.821,-587.69,0.0000,-1039.8,-1495.1,-734.11,-1142.9
1926.000000000,66.712,1521.3,1553.4,1193.0,224.05,2604.7,966.62,2.5546,5421.1,2758.1,3376.6,2110.9,0.0000,-5526.7,-6389.0,-876.14,-1713.7,-1229.2,-14705.,-86.913,-18476.,-5924.1,-3803.0,-2056.8,49.017,1746.2,1592.3,1205.8,245.64,2653.2,1686.6,0.0000,6414.2,4449.7,4252.8,3658.0,0.0000,-249.55,-75.865,-64.546,-32.678,-59.307,-587.69,0.0000,-1039.8,-1495.1,-734.08,-1142.8
1927.000000000,66.553,1517.0,1548.8,1185.3,223.38,2586.6,966.62,2.5549,5409.6,2758.2,3376.6,2111.0,0.0000,-5522.0,-6386.8,-873.84,-1712.9,-1224.8,-14703.,-86.888,-18474.,-5923.8,-3802.7,-2056.4,48.871,1741.0,1587.5,1197.9,244.83,2634.2,1686.6,0.0000,6402.7,4449.7,4252.8,3658.0,0.0000,-248.71,-75.609,-64.201,-32.581,-58.792,-587.69,0.0000,-1039.7,-1495.0,-734.06,-1142.7
1928.000000000,66.156,1512.6,1544.3,1177.6,222.70,2568.5,966.62,2.5552,5398.1,2758.2,3376.6,2111.1,0.0000,-5517.2,-6384.7,-871.54,-1712.1,-1220.5,-14702.,-86.864,-18472.,-5923.5,-3802.4,-2056.0,48.710,1735.3,1582.3,1189.7,243.95,2614.7,1686.6,0.0000,6390.9,4449.7,4252.8,3658.0,0.0000,-247.79,-75.330,-63.840,-32.473,-58.268,-587.69,0.0000,-1039.7,-1495.0,-734.04,-1142.6
1929.000000000,66.010,1508.0,1539.7,1170.0,221.95,2550.4,966.62,2.5555,5386.8,2758.2,3376.7,2111.2,0.0000,-5512.4,-6382.5,-869.23,-1711.3,-1216.1,-14701.,-86.839,-18470.,-5923.2,-3802.2,-2055.6,48.527,1728.7,1576.3,1181.1,242.97,2594.5,1686.6,0.0000,6378.6,4449.7,4252.8,3658.0,0.0000,-246.77,-75.017,-63.454,-32.351,-57.726,-587.69,0.0000,-1039.7,-1494.9,-734.02,-1142.5
1930.000000000,65.848,1503.2,1534.8,1162.3,221.17,2532.4,966.62,2.5765,5375.6,2758.3,3376.7,2111.2,0.0000,-5507.5,-6380.3,-866.92,-1710.5,-1211.6,-14699.,-86.815,-18468.,-5922.9,-3801.9,-2055.2,48.366,1723.0,1571.1,1173.2,242.09,2575.8,1686.6,0.0000,6367.3,4449.7,4252.8,3658.0,0.0000,-245.85,-74.739,-63.103,-32.244,-57.221,-587.69,0.0000,-1039.7,-1494.9,-733.99,-1142.4
1931.000000000,65.683,1498.8,1529.9,1154.7,220.44,2514.4,966.62,2.5854,5364.6,2758.3,3376.7,2111.3,0.0000,-5502.6,-6378.2,-864.61,-1709.7,-1207.2,-14698.,-86.791,-18466.,-5922.5,-3801.6,-2054.8,48.245,1718.7,1567.2,1165.9,241.41,2558.3,1686.6,0.0000,6356.7,4449.7,4252.8,3658.0,0.0000,-245.14,-74.521,-62.794,-32.163,-56.744,-587.69,0.0000,-1039.7,-1494.8,-733.97,-1142.3
1932.000000000,65.534,1494.6,1525.6,1147.2,219.80,2496.7,966.62,2.5857,5353.8,2758.4,3376.8,2111.4,0.0000,-5497.7,-6376.0,-862.29,-1708.9,-1202.7,-14696.,-86.766,-18464.,-5922.2,-3801.3,-2054.5,48.107,1713.8,1562.7,1158.4,240.65,2540.3,1686.6,0.0000,6345.8,4449.7,4252.8,3658.0,0.0000,-244.34,-74.279,-62.467,-32.071,-56.255,-587.69,0.0000,-1039.7,-1494.8,-733.95,-1142.2
1933.000000000,65.390,1490.3,1521.1,1139.6,219.08,2479.3,966.59,2.5860,5343.1,2758.4,3376.8,2111.5,0.0000,-5492.8,-6373.9,-859.97,-1708.1,-1198.3,-14695.,-86.742,-18462.,-5921.9,-3801.0,-2054.1,47.951,1708.2,1557.6,1150.5,239.80,2521.6,1686.6,0.0000,6334.4,4449.7,4252.8,3658.0,0.0000,-243.45,-74.008,-62.120,-31.967,-55.752,-587.69,0.0000,-1039.7,-1494.7,-733.92,-1142.1
1934.000000000,65.254,1485.9,1516.4,1132.3,218.34,2461.9,966.58,2.5863,5332.4,2758.5,3376.8,2111.6,0.0000,-5487.9,-6371.7,-857.65,-1707.3,-1193.8,-14693.,-86.718,-18460.,-5921.6,-3800.7,-2053.7,47.777,1702.0,1552.0,1142.4,238.86,2502.3,1686.6,0.0000,6322.7,4449.7,4252.8,3658.0,0.0000,-242.47,-73.710,-61.754,-31.851,-55.237,-587.69,0.0000,-1039.7,-1494.6,-733.90,-1142.0
1935.000000000,65.159,1481.3,1511.6,1125.1,217.60,2444.7,966.58,2.5866,5321.8,2758.5,3376.9,2111.7,0.0000,-5483.0,-6369.5,-855.32,-1706.5,-1189.3,-14692.,-86.693,-18457.,-5921.3,-3800.4,-2053.3,47.627,1696.7,1547.1,1134.7,238.04,2484.1,1686.6,0.0000,6311.7,4449.7,4252.8,3658.0,0.0000,-241.61,-73.447,-61.415,-31.751,-54.744,-587.69,0.0000,-1039.7,-1494.6,-733.88,-1141.9
1936.000000000,65.005,1476.7,1506.8,1117.8,216.89,2427.5,966.58,2.5869,5311.1,2758.6,3376.9,2111.8,0.0000,-5478.0,-6367.4,-852.98,-1705.7,-1184.8,-14690.,-86.669,-18455.,-5920.9,-3800.1,-2052.9,47.479,1691.4,1542.3,1127.1,237.23,2466.1,1686.6,0.0000,6300.7,4449.7,4252.8,3658.0,0.0000,-240.76,-73.190,-61.083,-31.653,-54.259,-587.69,0.0000,-1039.6,-1494.5,-733.85,-1141.8
1937.000000000,64.863,1472.1,1501.8,1110.4,216.17,2410.3,966.58,2.5872,5300.5,2758.6,3376.9,2111.9,0.0000,-5473.0,-6365.2,-850.64,-1704.8,-1180.2,-14689.,-86.645,-18453.,-5920.6,-3799.8,-2052.5,47.345,1686.6,1537.9,1119.9,236.49,2448.7,1686.6,0.0000,6290.2,4449.7,4252.8,3658.0,0.0000,-239.98,-72.956,-60.768,-31.563,-53.789,-587.69,0.0000,-1039.6,-1494.5,-733.83,-1141.7
1938.000000000,64.758,1467.7,1497.3,1103.2,215.49,2393.1,966.58,2.5875,5289.9,2758.7,3376.9,2112.0,0.0000,-5468.0,-6363.0,-848.31,-1704.0,-1175.6,-14687.,-86.620,-18451.,-5920.3,-3799.5,-2052.1,47.217,1682.1,1533.8,1112.8,235.78,2431.8,1686.6,0.0000,6279.9,4449.7,4252.8,3658.0,0.0000,-239.23,-72.732,-60.461,-31.478,-53.328,-587.69,0.0000,-1039.6,-1494.4,-733.81,-1141.6
1939.000000000,64.615,1463.6,1493.0,1096.0,214.84,2376.2,966.58,2.5878,5279.5,2758.7,3376.9,2112.1,0.0000,-5463.1,-6360.8,-845.97,-1703.2,-1171.1,-14686.,-86.596,-18449.,-5920.0,-3799.2,-2051.7,47.076,1677.1,1529.2,1105.5,235.01,2414.4,1686.6,0.0000,6269.4,4449.7,4252.8,3658.0,0.0000,-238.42,-72.489,-60.141,-31.384,-52.859,-587.69,0.0000,-1039.6,-1494.4,-733.78,-1141.5
1940.000000000,64.476,1459.4,1488.8,1088.9,214.16,2359.8,966.58,2.5881,5269.2,2758.5,3376.9,2112.2,0.0000,-5458.1,-6358.7,-843.63,-1702.4,-1166.5,-14684.,-86.572,-18447.,-5919.7,-3798.9,-2051.3,46.924,1671.6,1524.2,1098.0,234.18,2396.6,1686.6,0.0000,6258.6,4449.7,4252.8,3658.0,0.0000,-237.55,-72.228,-59.808,-31.282,-52.382,-587.69,0.0000,-1039.6,-1494.3,-733.76,-1141.4
1941.000000000,64.332,1455.1,1484.4,1081.9,213.46,2343.4,966.58,2.5884,5259.0,2758.5,3377.0,2112.3,0.0000,-5453.0,-6356.5,-841.29,-1701.6,-1161.9,-14683.,-86.548,-18445.,-5919.3,-3798.6,-2050.9,46.758,1665.7,1518.9,1090.3,233.29,2378.5,1686.6,0.0000,6247.6,4449.7,4252.8,3658.0,0.0000,-236.61,-71.947,-59.462,-31.172,-51.897,-587.69,0.0000,-1039.6,-1494.3,-733.74,-1141.3
1942.000000000,64.183,1451.4,1480.5,1074.9,212.86,2327.0,966.58,2.5887,5248.8,2758.6,3376.9,2112.4,0.0000,-5448.0,-6354.4,-838.95,-1700.8,-1157.3,-14681.,-86.524,-18442.,-5919.0,-3798.3,-2050.5,46.933,1669.2,1522.0,1086.6,233.67,2367.8,1686.6,0.0000,6241.1,4449.7,4252.8,3658.0,0.0000,-237.00,-72.069,-59.383,-31.236,-51.581,-587.69,0.0000,-1039.6,-1494.2,-733.71,-1141.2
1943.000000000,64.103,1449.4,1477.9,1068.1,212.62,2311.1,966.58,2.5890,5238.8,2758.6,3376.9,2112.5,0.0000,-5443.2,-6352.4,-836.63,-1700.0,-1152.7,-14680.,-86.500,-18440.,-5918.7,-3798.0,-2050.2,46.729,1664.7,1517.9,1079.6,232.98,2351.1,1686.6,0.0000,6231.0,4449.7,4252.8,3658.0,0.0000,-236.27,-71.851,-59.082,-31.152,-51.130,-587.69,0.0000,-1039.5,-1494.2,-733.69,-1141.1
1944.000000000,64.105,1446.8,1475.0,1061.5,212.06,2295.6,966.58,2.5893,5228.8,2758.7,3376.9,2112.6,0.0000,-5438.4,-6350.4,-834.31,-1699.2,-1148.1,-14678.,-86.476,-18438.,-5918.4,-3797.7,-2049.8,46.595,1659.9,1513.6,1072.5,232.24,2334.2,1686.6,0.0000,6220.8,4449.7,4252.8,3658.0,0.0000,-235.50,-71.621,-58.774,-31.063,-50.676,-587.69,0.0000,-1039.5,-1494.1,-733.67,-1141.0
1945.000000000,63.966,1443.5,1471.6,1055.3,211.49,2280.0,966.58,2.5927,5219.1,2758.7,3376.9,2112.7,0.0000,-5433.6,-6348.4,-831.99,-1698.4,-1143.5,-14677.,-86.452,-18436.,-5918.1,-3797.3,-2049.4,46.454,1654.9,1509.0,1065.4,231.47,2317.2,1686.6,0.0000,6210.5,4449.7,4252.8,3658.0,0.0000,-234.69,-71.379,-58.460,-30.969,-50.221,-587.69,0.0000,-1039.5,-1494.1,-733.64,-1140.9
1946.000000000,63.826,1439.7,1467.7,1048.9,211.01,2264.4,966.58,2.5954,5209.3,2758.8,3377.0,2112.8,0.0000,-5428.8,-6346.4,-829.67,-1697.6,-1138.8,-14675.,-86.428,-18434.,-5917.8,-3797.0,-2049.0,46.310,1649.8,1504.3,1058.2,230.69,2300.3,1686.6,0.0000,6200.2,4449.7,4252.8,3658.0,0.0000,-233.87,-71.133,-58.144,-30.873,-49.767,-587.69,0.0000,-1039.5,-1494.0,-733.62,-1140.8
1947.000000000,63.496,1435.6,1463.5,1042.5,210.39,2248.8,966.58,2.5957,5199.7,2758.8,3377.0,2112.9,0.0000,-5423.9,-6344.4,-827.35,-1696.8,-1134.2,-14674.,-86.404,-18431.,-5917.4,-3796.7,-2048.6,46.174,1644.9,1499.9,1051.3,229.95,2283.8,1686.6,0.0000,6190.2,4449.7,4252.8,3658.0,0.0000,-233.09,-70.899,-57.840,-30.783,-49.325,-587.69,0.0000,-1039.5,-1494.0,-733.60,-1140.7
1948.000000000,63.358,1431.6,1459.4,1035.9,209.65,2233.2,966.58,2.5960,5190.0,2758.9,3377.0,2112.9,0.0000,-5419.1,-6342.3,-825.02,-1696.0,-1129.5,-14672.,-86.380,-18429.,-5917.1,-3796.4,-2048.2,46.022,1639.5,1495.0,1044.1,229.12,2266.8,1686.6,0.0000,6179.9,4449.7,4252.8,3658.0,0.0000,-232.22,-70.640,-57.518,-30.681,-48.872,-587.69,0.0000,-1039.5,-1493.9,-733.57,-1140.6
1949.000000000,63.218,1427.6,1455.1,1029.3,208.98,2217.7,966.58,2.5963,5180.6,2758.9,3377.0,2113.0,0.0000,-5414.2,-6340.3,-822.71,-1695.2,-1124.9,-14670.,-86.356,-18427.,-5916.8,-3796.1,-2047.8,45.925,1636.1,1491.8,1037.8,228.57,2251.5,1686.6,0.0000,6170.6,4449.7,4252.8,3658.0,0.0000,-231.64,-70.467,-57.254,-30.617,-48.455,-587.69,0.0000,-1039.4,-1493.9,-733.55,-1140.6
1950.000000000,63.081,1430.3,1456.3,1023.0,209.19,2202.8,966.58,2.5966,5171.2,2759.0,3377.1,2113.2,0.0000,-5409.7,-6338.5,-820.46,-1694.4,-1120.2,-14669.,-86.334,-18425.,-5916.5,-3795.8,-2047.4,51.623,1699.2,1549.8,1055.8,237.25,2277.9,1686.6,1.0983,6186.5,4450.0,4253.1,3658.3,0.0000,-240.36,-73.154,-58.722,-31.783,-48.957,-587.69,-0.50149E-01,-1039.4,-1493.8,-733.53,-1140.5
1951.000000000,63.401,1448.9,1472.1,1017.9,212.59,2191.0,966.58,2.5969,5162.9,2759.0,3377.1,2113.3,0.0000,-5406.6,-6337.7,-818.36,-1693.8,-1115.6,-14667.,-86.313,-18423.,-5916.2,-3795.5,-2047.1,48.664,1739.6,1580.8,1059.3,242.08,2273.7,1686.6,0.0000,6183.7,4449.7,4252.8,3658.0,0.0000,-245.29,-74.636,-59.321,-32.446,-48.791,-587.69,0.0000,-1039.4,-1493.8,-733.51,-1140.4
1952.000000000,64.370,1470.2,1491.3,1015.3,214.94,2181.3,966.58,2.6002,5155.2,2759.1,3377.1,2113.4,0.0000,-5404.6,-6337.7,-816.29,-1693.4,-1111.1,-14666.,-86.291,-18420.,-5915.9,-3795.2,-2046.7,48.876,1741.2,1587.7,1054.0,242.89,2260.3,1686.6,0.0000,6175.3,4449.7,4252.8,3658.0,0.0000,-246.28,-74.953,-59.285,-32.587,-48.417,-587.69,0.0000,-1039.4,-1493.7,-733.48,-1140.3
1953.000000000,64.792,1483.9,1505.4,1015.1,216.28,2172.9,966.56,2.6261,5148.0,2759.1,3377.1,2113.5,0.0000,-5403.2,-6338.0,-814.25,-1693.0,-1106.7,-14664.,-86.269,-18418.,-5915.6,-3794.8,-2046.3,48.910,1742.4,1588.8,1048.4,242.62,2245.3,1686.6,0.0000,6166.2,4449.7,4252.8,3658.0,0.0000,-246.39,-74.998,-59.114,-32.608,-48.014,-587.69,0.0000,-1039.4,-1493.7,-733.46,-1140.2
1954.000000000,65.128,1490.6,1512.1,1013.8,218.14,2163.6,966.54,2.6265,5140.7,2759.2,3377.2,2113.6,0.0000,-5401.9,-6338.3,-812.26,-1692.6,-1102.4,-14662.,-86.246,-18416.,-5915.2,-3794.5,-2045.9,48.861,1740.6,1587.2,1042.3,242.17,2230.0,1686.6,0.0000,6156.9,4449.7,4252.8,3658.0,0.0000,-246.08,-74.915,-58.882,-32.574,-47.604,-587.69,0.0000,-1039.4,-1493.6,-733.44,-1140.1
1955.000000000,65.630,1492.8,1515.0,1011.7,219.13,2152.3,966.54,2.6267,5133.0,2759.2,3377.3,2113.7,0.0000,-5400.6,-6338.5,-810.26,-1692.1,-1098.0,-14661.,-86.222,-18414.,-5914.9,-3794.2,-2045.5,48.764,1737.2,1584.0,1035.9,241.58,2214.5,1686.6,0.0000,6147.5,4449.7,4252.8,3658.0,0.0000,-245.53,-74.759,-58.617,-32.509,-47.190,-587.69,0.0000,-1039.3,-1493.6,-733.41,-1140.0
1956.000000000,65.776,1492.8,1516.4,1008.1,219.08,2140.1,966.54,2.6309,5124.8,2759.3,3377.3,2113.7,0.0000,-5399.1,-6338.4,-808.23,-1691.7,-1093.5,-14659.,-86.199,-18412.,-5914.6,-3793.9,-2045.1,48.645,1733.0,1580.2,1029.4,240.91,2199.1,1686.6,0.0000,6138.2,4449.7,4252.8,3658.0,0.0000,-244.87,-74.568,-58.339,-32.430,-46.781,-587.69,0.0000,-1039.3,-1493.5,-733.39,-1139.9
1957.000000000,65.740,1491.9,1515.1,1003.6,218.71,2127.5,966.54,2.6327,5117.2,2759.3,3377.3,2113.8,0.0000,-5397.4,-6338.2,-806.25,-1691.1,-1089.0,-14658.,-86.175,-18409.,-5914.3,-3793.6,-2044.7,48.508,1728.1,1575.7,1022.9,240.17,2183.7,1686.6,0.0000,6128.8,4449.7,4252.8,3658.0,0.0000,-244.11,-74.349,-58.049,-32.339,-46.373,-587.69,0.0000,-1039.3,-1493.5,-733.37,-1139.8
1958.000000000,65.649,1489.8,1513.2,999.20,218.15,2113.9,966.54,2.6330,5109.7,2759.4,3377.4,2113.9,0.0000,-5395.5,-6337.8,-804.24,-1690.6,-1084.5,-14656.,-86.151,-18407.,-5914.0,-3793.2,-2044.4,48.360,1722.8,1570.9,1016.4,239.38,2168.4,1686.6,0.0000,6119.6,4449.7,4252.8,3658.0,0.0000,-243.31,-74.113,-57.753,-32.240,-45.968,-587.69,0.0000,-1039.3,-1493.4,-733.34,-1139.7
1959.000000000,65.528,1486.7,1511.6,994.05,217.47,2100.5,966.54,2.6333,5103.3,2759.8,3377.3,2114.0,0.0000,-5393.5,-6337.2,-802.18,-1690.0,-1079.9,-14654.,-86.127,-18405.,-5913.7,-3792.9,-2044.0,48.201,1717.1,1565.8,1009.8,238.54,2153.1,1686.6,0.0000,6110.3,4449.7,4252.8,3658.0,0.0000,-242.45,-73.859,-57.451,-32.134,-45.563,-587.69,0.0000,-1039.3,-1493.4,-733.32,-1139.6
1960.000000000,65.389,1483.8,1509.7,988.12,216.78,2088.8,966.54,2.6336,5098.3,2759.8,3377.3,2114.1,0.0000,-5391.3,-6336.6,-800.09,-1689.4,-1075.4,-14653.,-86.103,-18403.,-5913.3,-3792.6,-2043.6,48.031,1711.1,1560.2,1003.1,237.64,2137.7,1686.6,0.0000,6101.0,4449.7,4252.8,3658.0,0.0000,-241.53,-73.586,-57.139,-32.021,-45.157,-587.69,0.0000,-1039.3,-1493.3,-733.30,-1139.5
1961.000000000,65.236,1481.3,1507.3,982.15,216.05,2078.0,966.54,2.6338,5092.6,2759.6,3377.3,2114.1,0.0000,-5389.0,-6335.8,-797.98,-1688.8,-1070.8,-14651.,-86.079,-18401.,-5913.0,-3792.3,-2043.2,47.871,1705.4,1555.0,996.73,236.80,2122.9,1686.6,0.0000,6092.0,4449.7,4252.8,3658.0,0.0000,-240.65,-73.327,-56.841,-31.914,-44.764,-587.69,0.0000,-1039.2,-1493.3,-733.27,-1139.4
1962.000000000,65.076,1477.4,1503.2,977.01,215.31,2067.6,966.54,2.6597,5086.2,2759.6,3377.3,2114.3,0.0000,-5386.4,-6334.9,-795.86,-1688.2,-1066.2,-14650.,-86.055,-18398.,-5912.7,-3792.0,-2042.8,47.699,1699.3,1549.4,990.20,235.90,2107.8,1686.6,0.0000,6082.9,4449.7,4252.8,3658.0,0.0000,-239.73,-73.051,-56.533,-31.800,-44.367,-587.69,0.0000,-1039.2,-1493.2,-733.25,-1139.3
1963.000000000,64.879,1473.1,1498.1,971.62,214.50,2055.3,966.54,2.6619,5079.1,2759.7,3377.3,2114.4,0.0000,-5383.6,-6333.9,-793.73,-1687.5,-1061.6,-14648.,-86.032,-18396.,-5912.4,-3791.6,-2042.4,47.523,1693.0,1543.7,983.64,234.98,2092.8,1686.6,0.0000,6073.8,4449.7,4252.8,3658.0,0.0000,-238.77,-72.765,-56.222,-31.682,-43.971,-587.69,0.0000,-1039.2,-1493.2,-733.23,-1139.2
1964.000000000,64.679,1469.6,1493.3,966.33,213.71,2042.4,966.54,2.6648,5071.3,2759.7,3377.3,2114.5,0.0000,-5380.6,-6332.8,-791.59,-1686.9,-1056.9,-14646.,-86.008,-18394.,-5912.1,-3791.3,-2042.0,47.341,1686.5,1537.8,977.16,234.03,2078.0,1686.6,0.0000,6064.8,4449.7,4252.8,3658.0,0.0000,-237.79,-72.472,-55.911,-31.561,-43.581,-587.69,0.0000,-1039.2,-1493.1,-733.20,-1139.1
1965.000000000,64.505,1465.9,1489.1,960.76,212.93,2028.6,966.54,2.6768,5063.3,2759.8,3377.4,2114.6,0.0000,-5377.4,-6331.7,-789.44,-1686.2,-1052.3,-14645.,-85.984,-18392.,-5911.8,-3791.0,-2041.7,47.164,1680.2,1532.0,970.67,233.11,2063.1,1686.6,0.0000,6055.8,4449.7,4252.8,3658.0,0.0000,-236.82,-72.184,-55.602,-31.442,-43.191,-587.69,0.0000,-1039.2,-1493.1,-733.18,-1139.1
1966.000000000,64.288,1461.2,1484.9,954.86,212.17,2014.7,966.53,2.6771,5055.0,2759.8,3377.4,2114.7,0.0000,-5374.1,-6330.5,-787.30,-1685.6,-1047.6,-14643.,-85.960,-18390.,-5911.5,-3790.7,-2041.3,47.043,1675.9,1528.1,965.62,232.47,2051.4,1686.6,0.0000,6048.7,4449.7,4252.8,3658.0,0.0000,-236.14,-71.983,-55.368,-31.362,-42.869,-587.69,0.0000,-1039.2,-1493.0,-733.16,-1139.0
1967.000000000,64.101,1463.7,1486.1,949.08,212.39,2002.0,966.52,2.6774,5046.6,2759.9,3377.4,2114.8,0.0000,-5371.1,-6329.5,-785.23,-1685.0,-1043.0,-14641.,-85.939,-18387.,-5911.1,-3790.3,-2040.9,122.42,1782.1,1641.6,988.27,244.24,2084.8,1686.6,15.928,6069.8,4452.5,4255.6,3660.8,0.0000,-245.06,-75.881,-56.909,-32.567,-43.470,-587.69,-0.72727,-1039.2,-1493.0,-733.15,-1138.9
1968.000000000,64.452,1482.7,1501.8,944.14,215.77,1991.9,966.51,2.6777,5039.1,2759.9,3377.4,2114.9,0.0000,-5369.4,-6329.4,-783.29,-1684.5,-1038.5,-14640.,-85.918,-18385.,-5910.8,-3790.0,-2040.5,49.608,1767.2,1611.4,986.43,244.88,2075.6,1686.6,0.0000,6063.4,4450.0,4253.4,3658.2,0.0000,-248.90,-75.891,-57.338,-33.074,-43.240,-587.69,0.0000,-1039.1,-1492.9,-733.11,-1138.8
1969.000000000,65.390,1501.8,1520.3,941.98,217.62,1983.7,966.48,2.6780,5032.4,2759.9,3377.4,2115.0,0.0000,-5368.8,-6330.1,-781.37,-1684.2,-1034.0,-14638.,-85.896,-18383.,-5910.5,-3789.7,-2040.1,49.720,1771.3,1615.1,981.51,245.10,2062.2,1686.6,0.0000,6054.9,4449.8,4253.0,3658.0,0.0000,-249.42,-76.061,-57.243,-33.147,-42.888,-587.69,0.0000,-1039.1,-1492.9,-733.09,-1138.7
1970.000000000,65.685,1512.7,1531.8,942.10,218.77,1976.9,966.48,2.6783,5026.0,2760.0,3377.5,2115.1,0.0000,-5368.5,-6331.0,-779.48,-1683.9,-1029.7,-14636.,-85.874,-18381.,-5910.2,-3789.4,-2039.7,49.693,1770.3,1614.2,976.04,244.82,2048.5,1686.6,0.0000,6046.4,4449.7,4252.8,3658.0,0.0000,-249.25,-76.019,-57.050,-33.129,-42.529,-587.69,0.0000,-1039.1,-1492.8,-733.06,-1138.6
1971.000000000,66.009,1518.0,1536.3,940.86,220.43,1969.1,966.48,2.6785,5019.8,2760.0,3377.5,2115.2,0.0000,-5368.2,-6331.7,-777.61,-1683.6,-1025.4,-14635.,-85.851,-18379.,-5909.9,-3789.0,-2039.4,49.598,1766.9,1611.1,970.31,244.28,2034.7,1686.6,0.0000,6038.0,4449.7,4252.8,3658.0,0.0000,-248.73,-75.871,-56.810,-33.065,-42.168,-587.69,0.0000,-1039.1,-1492.8,-733.04,-1138.5
1972.000000000,66.415,1518.5,1537.6,938.66,221.01,1959.6,966.48,2.6788,5012.9,2760.1,3377.5,2115.2,0.0000,-5367.9,-6332.2,-775.75,-1683.2,-1021.1,-14633.,-85.827,-18376.,-5909.6,-3788.7,-2039.0,49.459,1761.9,1606.6,964.33,243.53,2020.8,1686.6,0.0000,6029.6,4449.7,4252.8,3658.0,0.0000,-248.00,-75.656,-56.539,-32.973,-41.804,-587.69,0.0000,-1039.0,-1492.7,-733.02,-1138.4
1973.000000000,66.465,1517.0,1537.5,935.77,220.68,1948.8,966.48,2.6791,5005.9,2760.1,3377.5,2115.3,0.0000,-5367.3,-6332.4,-773.86,-1682.8,-1016.7,-14631.,-85.804,-18374.,-5909.3,-3788.4,-2038.6,49.290,1755.9,1601.1,958.13,242.65,2006.6,1686.6,0.0000,6021.0,4449.7,4252.8,3658.0,0.0000,-247.11,-75.393,-56.244,-32.860,-41.436,-587.69,0.0000,-1039.0,-1492.7,-732.99,-1138.3
1974.000000000,66.371,1514.6,1534.7,931.65,220.07,1937.7,966.48,2.6794,4998.9,2760.2,3377.5,2115.4,0.0000,-5366.4,-6332.5,-771.97,-1682.3,-1012.3,-14630.,-85.781,-18372.,-5909.0,-3788.0,-2038.2,49.105,1749.4,1595.1,951.89,241.70,1992.4,1686.6,0.0000,6012.4,4449.7,4252.8,3658.0,0.0000,-246.15,-75.106,-55.941,-32.737,-41.070,-587.69,0.0000,-1039.0,-1492.6,-732.97,-1138.2
1975.000000000,66.229,1511.1,1531.4,927.84,219.34,1926.0,966.48,2.6796,4993.0,2760.2,3377.6,2115.5,0.0000,-5365.2,-6332.3,-770.09,-1681.9,-1007.8,-14628.,-85.757,-18370.,-5908.6,-3787.7,-2037.8,48.916,1742.6,1589.0,945.70,240.72,1978.5,1686.6,0.0000,6004.0,4449.7,4252.8,3658.0,0.0000,-245.16,-74.810,-55.636,-32.610,-40.709,-587.69,0.0000,-1039.0,-1492.6,-732.95,-1138.1
1976.000000000,66.062,1506.8,1528.4,923.53,218.51,1913.9,966.48,2.6799,4986.4,2760.3,3377.6,2115.5,0.0000,-5363.8,-6332.0,-768.17,-1681.3,-1003.4,-14626.,-85.733,-18368.,-5908.3,-3787.4,-2037.4,48.721,1735.7,1582.6,939.55,239.72,1964.7,1686.6,0.0000,5995.6,4449.7,4252.8,3658.0,0.0000,-244.15,-74.505,-55.331,-32.481,-40.352,-587.69,0.0000,-1039.0,-1492.5,-732.92,-1138.0
1977.000000000,65.904,1503.4,1525.5,918.22,217.66,1902.9,966.48,2.6802,4981.5,2760.3,3377.6,2115.6,0.0000,-5362.2,-6331.5,-766.21,-1680.8,-998.88,-14625.,-85.710,-18365.,-5908.0,-3787.0,-2037.1,48.521,1728.5,1576.1,933.38,238.70,1950.9,1686.6,0.0000,5987.3,4449.7,4252.8,3658.0,0.0000,-243.10,-74.189,-55.021,-32.347,-39.996,-587.69,0.0000,-1038.9,-1492.5,-732.90,-1137.9
1978.000000000,65.791,1499.5,1521.4,913.32,216.80,1893.2,966.49,2.6805,4977.4,2760.4,3377.7,2115.7,0.0000,-5360.3,-6330.8,-764.22,-1680.2,-994.38,-14623.,-85.686,-18363.,-5907.7,-3786.7,-2036.7,48.350,1722.5,1570.6,927.79,237.82,1938.3,1686.6,0.0000,5979.7,4449.7,4252.8,3658.0,0.0000,-242.20,-73.917,-54.746,-32.234,-39.665,-587.69,0.0000,-1038.9,-1492.4,-732.87,-1137.8
1979.000000000,65.602,1494.6,1516.8,908.64,215.91,1883.6,966.49,2.6807,4972.1,2760.6,3377.7,2115.8,0.0000,-5358.3,-6330.0,-762.23,-1679.6,-989.86,-14621.,-85.663,-18361.,-5907.4,-3786.4,-2036.3,48.173,1716.1,1564.8,922.13,236.91,1925.6,1686.6,0.0000,5972.0,4449.7,4252.8,3658.0,0.0000,-241.26,-73.633,-54.465,-32.115,-39.333,-587.69,0.0000,-1038.9,-1492.4,-732.85,-1137.8
1980.000000000,65.473,1489.9,1512.3,903.56,215.08,1874.7,966.49,2.6810,4966.5,2760.8,3377.7,2115.9,0.0000,-5356.0,-6329.1,-760.23,-1679.0,-985.33,-14620.,-85.639,-18359.,-5907.1,-3786.0,-2035.9,47.987,1709.5,1558.8,916.38,235.95,1912.8,1686.6,0.0000,5964.2,4449.7,4252.8,3658.0,0.0000,-240.28,-73.335,-54.176,-31.991,-38.999,-587.69,0.0000,-1038.9,-1492.3,-732.83,-1137.7
1981.000000000,65.377,1486.6,1508.6,898.36,214.27,1863.7,966.48,2.6813,4960.4,2760.9,3377.7,2115.9,0.0000,-5353.6,-6328.1,-758.23,-1678.4,-980.79,-14618.,-85.616,-18357.,-5906.7,-3785.7,-2035.5,47.849,1704.6,1554.3,911.26,235.23,1901.0,1686.6,0.0000,5957.1,4449.7,4252.8,3658.0,0.0000,-239.53,-73.110,-53.933,-31.899,-38.689,-587.69,0.0000,-1038.9,-1492.3,-732.80,-1137.6
1982.000000000,65.203,1482.7,1505.0,893.41,213.58,1852.2,966.44,2.6815,4953.7,2761.0,3377.7,2116.0,0.0000,-5351.0,-6327.1,-756.23,-1677.8,-976.25,-14616.,-85.592,-18354.,-5906.4,-3785.4,-2035.1,47.678,1698.5,1548.8,905.85,234.36,1888.9,1686.6,0.0000,5949.7,4449.7,4252.8,3658.0,0.0000,-238.63,-72.836,-53.664,-31.786,-38.371,-587.69,0.0000,-1038.8,-1492.2,-732.78,-1137.5
1983.000000000,65.044,1478.0,1500.6,888.48,212.81,1840.4,966.44,2.6818,4946.9,2761.0,3377.7,2116.1,0.0000,-5348.3,-6326.0,-754.22,-1677.2,-971.70,-14615.,-85.569,-18352.,-5906.1,-3785.0,-2034.7,47.493,1691.9,1542.8,900.23,233.41,1876.4,1686.6,0.0000,5942.2,4449.7,4252.8,3658.0,0.0000,-237.65,-72.539,-53.381,-31.662,-38.046,-587.69,0.0000,-1038.8,-1492.2,-732.76,-1137.4
1984.000000000,64.866,1473.3,1495.9,883.55,212.02,1828.6,966.45,2.6821,4939.6,2761.0,3377.8,2116.2,0.0000,-5345.5,-6324.9,-752.21,-1676.6,-967.15,-14613.,-85.546,-18350.,-5905.8,-3784.7,-2034.4,47.309,1685.4,1536.8,894.66,232.47,1864.0,1686.6,0.0000,5934.7,4449.7,4252.8,3658.0,0.0000,-236.67,-72.241,-53.099,-31.539,-37.724,-587.69,0.0000,-1038.8,-1492.1,-732.73,-1137.3
1985.000000000,64.688,1468.6,1492.1,878.70,211.25,1816.9,966.45,2.6823,4932.5,2761.1,3377.8,2116.3,0.0000,-5342.6,-6323.7,-750.20,-1675.9,-962.61,-14611.,-85.522,-18348.,-5905.5,-3784.4,-2034.0,47.132,1679.1,1531.0,889.23,231.57,1851.9,1686.6,0.0000,5927.4,4449.7,4252.8,3658.0,0.0000,-235.73,-71.955,-52.826,-31.422,-37.435,-587.69,0.0000,-1038.8,-1492.1,-732.71,-1137.2
1986.000000000,64.515,1463.3,1488.4,873.54,210.47,1805.4,966.44,2.6826,4925.2,2761.1,3377.8,2116.4,0.0000,-5339.7,-6322.4,-748.19,-1675.3,-958.09,-14610.,-85.499,-18346.,-5905.2,-3784.0,-2033.6,46.962,1673.0,1525.5,883.95,230.70,1840.1,1686.6,0.0000,5920.2,4449.7,4252.8,3658.0,0.0000,-234.82,-71.679,-52.562,-31.308,-37.152,-587.69,0.0000,-1038.8,-1492.0,-732.69,-1137.1
1987.000000000,64.410,1458.5,1483.5,868.38,209.69,1794.1,966.42,2.6829,4918.1,2761.2,3377.8,2116.4,0.0000,-5336.7,-6321.0,-746.17,-1674.6,-953.56,-14608.,-85.475,-18343.,-5904.9,-3783.7,-2033.2,46.792,1666.9,1520.0,878.68,229.83,1828.3,1686.6,0.0000,5913.1,4449.7,4252.8,3658.0,0.0000,-233.91,-71.401,-52.297,-31.195,-36.871,-587.69,0.0000,-1038.7,-1492.0,-732.66,-1137.0
1988.000000000,64.243,1453.9,1478.4,863.23,208.91,1782.8,966.42,2.6831,4911.3,2761.2,3377.8,2116.6,0.0000,-5333.6,-6319.6,-744.16,-1673.9,-949.04,-14606.,-85.452,-18341.,-5904.5,-3783.3,-2032.8,46.623,1660.9,1514.5,873.48,228.96,1816.7,1686.6,0.0000,5906.1,4449.7,4252.8,3658.0,0.0000,-233.00,-71.125,-52.036,-31.082,-36.593,-587.69,0.0000,-1038.7,-1491.9,-732.64,-1136.9
1989.000000000,64.068,1448.8,1473.2,858.07,208.12,1772.2,966.42,2.6834,4904.4,2761.3,3377.9,2116.7,0.0000,-5330.3,-6318.1,-742.15,-1673.2,-944.51,-14604.,-85.429,-18339.,-5904.2,-3783.0,-2032.4,46.449,1654.7,1508.8,868.20,228.07,1805.0,1686.6,0.0000,5899.0,4449.7,4252.8,3658.0,0.0000,-232.07,-70.841,-51.769,-30.966,-36.312,-587.69,0.0000,-1038.7,-1491.9,-732.62,-1136.8
1990.000000000,63.896,1443.6,1467.7,853.09,207.35,1761.2,966.42,2.6837,4897.4,2761.3,3377.9,2116.8,0.0000,-5326.9,-6316.6,-740.14,-1672.5,-939.97,-14603.,-85.405,-18337.,-5903.9,-3782.7,-2032.1,46.281,1648.7,1503.4,863.03,227.21,1793.4,1686.6,0.0000,5892.0,4449.7,4252.8,3658.0,0.0000,-231.17,-70.566,-51.510,-30.854,-36.037,-587.69,0.0000,-1038.7,-1491.8,-732.59,-1136.7
1991.000000000,63.678,1438.6,1462.5,848.39,206.61,1750.3,966.42,2.6839,4890.4,2761.4,3377.9,2116.9,0.0000,-5323.4,-6315.0,-738.13,-1671.8,-935.43,-14601.,-85.382,-18335.,-5903.6,-3782.3,-2031.7,46.119,1643.0,1498.1,857.98,226.38,1782.1,1686.6,0.0000,5885.2,4449.7,4252.8,3658.0,0.0000,-230.29,-70.300,-51.257,-30.746,-35.767,-587.69,0.0000,-1038.7,-1491.8,-732.57,-1136.6
1992.000000000,63.492,1433.6,1457.3,843.81,205.87,1739.3,966.41,2.6842,4883.7,2761.5,3377.9,2117.0,0.0000,-5319.9,-6313.3,-736.12,-1671.1,-930.88,-14599.,-85.359,-18332.,-5903.3,-3782.0,-2031.3,45.958,1637.2,1492.9,852.97,225.56,1770.9,1686.6,0.0000,5878.4,4449.7,4252.8,3658.0,0.0000,-229.43,-70.035,-51.007,-30.638,-35.499,-587.69,0.0000,-1038.6,-1491.7,-732.54,-1136.5
1993.000000000,63.327,1429.0,1452.2,839.00,205.14,1728.3,966.38,2.6819,4877.1,2761.8,3377.9,2117.0,0.0000,-5316.2,-6311.7,-734.12,-1670.4,-926.33,-14598.,-85.335,-18330.,-5903.0,-3781.6,-2030.9,45.797,1631.5,1487.6,847.98,224.73,1759.8,1686.6,0.0000,5871.6,4449.7,4252.8,3658.0,0.0000,-228.56,-69.770,-50.757,-30.531,-35.233,-587.69,0.0000,-1038.6,-1491.7,-732.52,-1136.4
1994.000000000,63.162,1424.3,1447.1,834.46,204.41,1717.6,966.38,2.6799,4870.6,2761.9,3377.9,2117.1,0.0000,-5312.4,-6309.9,-732.12,-1669.7,-921.78,-14596.,-85.312,-18328.,-5902.7,-3781.3,-2030.5,45.638,1625.8,1482.5,843.05,223.92,1748.8,1686.6,0.0000,5865.0,4449.7,4252.8,3658.0,0.0000,-227.70,-69.508,-50.510,-30.425,-34.970,-587.69,0.0000,-1038.6,-1491.6,-732.50,-1136.4
1995.000000000,62.999,1419.5,1442.3,829.99,203.70,1707.0,966.38,2.6802,4864.0,2761.9,3378.0,2117.2,0.0000,-5308.6,-6308.2,-730.13,-1668.9,-917.23,-14594.,-85.289,-18326.,-5902.3,-3781.0,-2030.1,45.488,1620.5,1477.6,838.18,223.15,1737.8,1686.6,0.0000,5858.3,4449.7,4252.8,3658.0,0.0000,-226.88,-69.259,-50.270,-30.326,-34.709,-587.69,0.0000,-1038.6,-1491.6,-732.47,-1136.3
1996.000000000,62.841,1414.6,1437.5,825.26,203.02,1696.4,966.38,2.6805,4857.8,2762.0,3378.0,2117.3,0.0000,-5304.7,-6306.4,-728.14,-1668.2,-912.68,-14593.,-85.266,-18324.,-5902.0,-3780.6,-2029.8,45.360,1615.9,1473.5,834.11,222.49,1728.7,1686.6,0.0000,5852.8,4449.7,4252.8,3658.0,0.0000,-226.17,-69.043,-50.066,-30.240,-34.486,-587.69,0.0000,-1038.6,-1491.5,-732.45,-1136.2
1997.000000000,62.691,1410.3,1434.4,820.62,202.38,1685.7,966.38,2.6807,4851.3,2762.0,3378.1,2117.4,0.0000,-5300.9,-6304.6,-726.17,-1667.5,-908.13,-14591.,-85.242,-18321.,-5901.7,-3780.3,-2029.4,45.210,1610.6,1468.6,829.35,221.72,1718.0,1686.6,0.0000,5846.3,4449.7,4252.8,3658.0,0.0000,-225.35,-68.792,-49.829,-30.140,-34.231,-587.69,0.0000,-1038.5,-1491.5,-732.43,-1136.1
1998.000000000,62.547,1406.2,1430.0,816.05,201.73,1675.4,966.38,2.6810,4844.9,2762.1,3378.2,2117.4,0.0000,-5297.0,-6302.8,-724.20,-1666.7,-903.58,-14589.,-85.219,-18319.,-5901.4,-3779.9,-2029.0,45.061,1605.3,1463.8,824.65,220.96,1707.5,1686.6,0.0000,5840.0,4449.7,4252.8,3658.0,0.0000,-224.55,-68.546,-49.595,-30.041,-33.979,-587.69,0.0000,-1038.5,-1491.4,-732.40,-1136.0
1999.000000000,62.447,1401.8,1425.5,811.51,201.09,1665.4,966.38,2.6812,4838.7,2762.1,3378.2,2117.5,0.0000,-5293.1,-6300.9,-722.25,-1666.0,-899.03,-14587.,-85.196,-18317.,-5901.1,-3779.6,-2028.6,44.927,1600.5,1459.4,820.22,220.26,1697.5,1686.6,0.0000,5833.9,4449.7,4252.8,3658.0,0.0000,-223.81,-68.320,-49.378,-29.951,-33.739,-587.69,0.0000,-1038.5,-1491.4,-732.38,-1135.9
2000.000000000,62.351,1397.4,1421.0,806.96,200.47,1655.5,966.38,2.6815,4832.7,2762.2,3378.3,2117.6,0.0000,-5289.1,-6299.1,-720.30,-1665.2,-894.48,-14586.,-85.173,-18315.,-5900.8,-3779.2,-2028.2,44.770,1594.9,1454.3,815.43,219.46,1686.8,1686.6,0.0000,5827.4,4449.7,4252.8,3658.0,0.0000,-222.96,-68.060,-49.137,-29.847,-33.486,-587.69,0.0000,-1038.5,-1491.3,-732.36,-1135.8
2001.000000000,62.211,1392.9,1417.0,802.89,199.76,1645.3,966.38,2.6817,4826.6,2762.2,3378.3,2117.7,0.0000,-5285.1,-6297.2,-718.36,-1664.5,-889.93,-14584.,-85.150,-18312.,-5900.5,-3778.9,-2027.9,44.608,1589.1,1449.0,810.55,218.63,1676.0,1686.6,0.0000,5820.9,4449.7,4252.8,3658.0,0.0000,-222.08,-67.791,-48.890,-29.738,-33.229,-587.69,0.0000,-1038.4,-1491.3,-732.33,-1135.7
2002.000000000,62.046,1388.4,1412.9,798.54,199.05,1635.1,966.38,2.6820,4820.8,2762.3,3378.3,2117.8,0.0000,-5281.1,-6295.3,-716.43,-1663.7,-885.36,-14582.,-85.127,-18310.,-5900.2,-3778.6,-2027.5,44.450,1583.5,1443.9,805.78,217.83,1665.3,1686.6,0.0000,5814.5,4449.7,4252.8,3658.0,0.0000,-221.22,-67.530,-48.650,-29.633,-32.977,-587.69,0.0000,-1038.4,-1491.2,-732.31,-1135.6
2003.000000000,61.890,1383.8,1408.4,794.15,198.35,1625.2,966.38,2.6823,4814.7,2762.3,3378.3,2117.9,0.0000,-5277.0,-6293.4,-714.51,-1662.9,-880.80,-14580.,-85.104,-18308.,-5899.8,-3778.2,-2027.1,44.302,1578.2,1439.1,801.17,217.07,1655.0,1686.6,0.0000,5808.2,4449.7,4252.8,3658.0,0.0000,-220.41,-67.283,-48.420,-29.535,-32.733,-587.69,0.0000,-1038.4,-1491.2,-732.28,-1135.5
2004.000000000,61.772,1379.2,1403.9,789.70,197.68,1615.5,966.38,2.6825,4808.8,2762.4,3378.3,2118.0,0.0000,-5272.9,-6291.5,-712.60,-1662.2,-876.23,-14579.,-85.081,-18306.,-5899.5,-3777.9,-2026.7,44.153,1572.9,1434.2,796.56,216.31,1644.7,1686.6,0.0000,5802.0,4449.7,4252.8,3658.0,0.0000,-219.60,-67.034,-48.189,-29.435,-32.488,-587.69,0.0000,-1038.4,-1491.1,-732.26,-1135.4
2005.000000000,61.771,1374.7,1399.3,785.28,197.00,1605.7,966.38,2.6828,4803.0,2762.4,3378.3,2118.0,0.0000,-5268.8,-6289.5,-710.71,-1661.4,-871.67,-14577.,-85.057,-18303.,-5899.2,-3777.5,-2026.3,44.003,1567.6,1429.4,791.96,215.54,1634.5,1686.6,0.0000,5795.8,4449.7,4252.8,3658.0,0.0000,-218.78,-66.785,-47.958,-29.336,-32.245,-587.69,0.0000,-1038.4,-1491.1,-732.24,-1135.3
2006.000000000,61.625,1370.2,1394.8,780.90,196.33,1595.8,966.38,2.6830,4797.0,2762.5,3378.4,2118.1,0.0000,-5264.5,-6287.6,-708.82,-1660.6,-867.11,-14575.,-85.034,-18301.,-5898.9,-3777.2,-2026.0,43.856,1562.3,1424.6,787.41,214.79,1624.3,1686.6,0.0000,5789.6,4449.7,4252.8,3658.0,0.0000,-217.98,-66.539,-47.731,-29.237,-32.004,-587.69,0.0000,-1038.3,-1491.0,-732.21,-1135.2
2007.000000000,61.520,1365.9,1390.3,776.54,195.71,1585.9,966.38,2.6833,4791.0,2762.5,3378.4,2118.3,0.0000,-5260.3,-6285.6,-706.95,-1659.8,-862.55,-14574.,-85.011,-18299.,-5898.6,-3776.8,-2025.6,43.755,1558.8,1421.3,783.71,214.26,1615.8,1686.6,0.0000,5784.5,4449.7,4252.8,3658.0,0.0000,-217.40,-66.364,-47.554,-29.170,-31.798,-587.69,0.0000,-1038.3,-1491.0,-732.19,-1135.1
2008.000000000,61.380,1361.9,1386.1,772.23,195.18,1576.3,966.38,2.5165,4785.0,2762.6,3378.4,2118.4,0.0000,-5256.0,-6283.7,-705.10,-1659.0,-857.97,-14572.,-84.988,-18297.,-5898.3,-3776.5,-2025.2,43.628,1554.2,1417.2,779.50,213.60,1606.3,1686.6,0.0000,5778.8,4449.7,4252.8,3658.0,0.0000,-216.70,-66.149,-47.348,-29.085,-31.572,-587.69,0.0000,-1038.3,-1490.9,-732.17,-1135.0
2009.000000000,61.216,1358.3,1382.2,767.99,194.59,1566.9,966.38,2.4111,4779.3,2762.6,3378.5,2118.5,0.0000,-5251.7,-6281.7,-703.26,-1658.2,-853.40,-14570.,-84.966,-18294.,-5898.0,-3776.1,-2024.8,43.497,1549.6,1412.9,775.26,212.93,1596.8,1686.6,0.0000,5773.0,4449.7,4252.8,3658.0,0.0000,-215.97,-65.928,-47.138,-28.998,-31.345,-587.69,0.0000,-1038.3,-1490.9,-732.14,-1134.9
2010.000000000,61.014,1354.4,1378.2,763.84,193.99,1557.7,966.38,2.4113,4773.4,2762.7,3378.5,2118.6,0.0000,-5247.4,-6279.8,-701.44,-1657.5,-848.82,-14568.,-84.943,-18292.,-5897.7,-3775.8,-2024.4,43.368,1545.0,1408.8,771.06,212.27,1587.3,1686.6,0.0000,5767.3,4449.7,4252.8,3658.0,0.0000,-215.26,-65.711,-46.931,-28.912,-31.120,-587.69,0.0000,-1038.2,-1490.8,-732.12,-1134.9
2011.000000000,60.880,1350.5,1374.1,759.87,193.37,1548.6,966.39,2.4116,4767.7,2762.7,3378.5,2118.7,0.0000,-5243.0,-6277.8,-699.64,-1656.7,-844.24,-14567.,-84.920,-18290.,-5897.4,-3775.5,-2024.0,43.238,1540.3,1404.5,766.86,211.60,1577.9,1686.6,0.0000,5761.5,4449.7,4252.8,3658.0,0.0000,-214.54,-65.492,-46.724,-28.825,-30.896,-587.69,0.0000,-1038.2,-1490.8,-732.09,-1134.8
2012.000000000,60.733,1346.8,1370.1,755.80,192.82,1539.5,966.39,2.4118,4762.0,2762.8,3378.6,2118.8,0.0000,-5238.7,-6275.9,-697.86,-1655.9,-839.67,-14565.,-84.897,-18288.,-5897.0,-3775.1,-2023.7,43.187,1538.5,1402.9,764.29,211.32,1571.8,1686.6,0.0000,5757.8,4449.7,4252.8,3658.0,0.0000,-214.21,-65.392,-46.609,-28.791,-30.741,-587.69,0.0000,-1038.2,-1490.7,-732.07,-1134.7
2013.000000000,60.578,1343.9,1366.8,751.81,192.44,1530.6,966.39,2.4120,4756.4,2762.8,3378.6,2118.9,0.0000,-5234.4,-6274.0,-696.11,-1655.1,-835.09,-14563.,-84.874,-18285.,-5896.7,-3774.8,-2023.3,43.192,1538.7,1403.0,762.54,211.31,1567.2,1686.6,0.10839,5755.1,4449.7,4252.9,3658.1,0.0000,-214.16,-65.378,-46.549,-28.794,-30.615,-587.69,-0.49490E-02,-1038.2,-1490.7,-732.05,-1134.6
2014.000000000,60.508,1342.7,1365.2,748.02,192.25,1522.2,966.39,2.4123,4750.8,2762.8,3378.6,2119.0,0.0000,-5230.3,-6272.2,-694.41,-1654.3,-830.52,-14561.,-84.853,-18283.,-5896.4,-3774.4,-2022.9,43.476,1546.5,1410.0,766.22,212.52,1573.7,1686.6,1.9021,5759.5,4450.8,4255.5,3661.1,0.0000,-215.02,-65.660,-46.729,-28.921,-30.701,-587.69,-0.86849E-01,-1038.2,-1490.6,-732.04,-1134.5
2015.000000000,60.499,1345.5,1367.1,744.74,192.62,1514.6,966.39,2.4125,4745.5,2762.9,3378.6,2119.0,0.0000,-5226.5,-6270.7,-692.78,-1653.6,-825.99,-14560.,-84.832,-18281.,-5896.1,-3774.1,-2022.5,45.306,1582.0,1449.2,784.69,223.27,1593.5,1686.6,8.4035,5771.5,4454.0,4260.8,3663.8,0.0000,-218.32,-67.032,-47.288,-29.418,-30.915,-587.69,-0.38369,-1038.2,-1490.6,-732.04,-1134.4
2016.000000000,60.692,1353.6,1373.9,742.37,194.00,1508.3,966.39,2.4127,4740.8,2763.0,3378.7,2119.1,0.0000,-5223.3,-6269.6,-691.22,-1652.9,-821.51,-14558.,-84.812,-18279.,-5895.8,-3773.7,-2022.2,44.450,1583.5,1443.9,773.26,217.27,1595.9,1686.6,0.0000,5763.8,4449.7,4263.3,3659.7,0.0000,-220.20,-67.229,-47.524,-29.633,-30.870,-587.69,0.0000,-1038.1,-1490.6,-732.03,-1134.3
2017.000000000,61.233,1364.2,1383.1,741.11,195.33,1502.9,966.39,2.4130,4736.3,2763.0,3378.7,2119.3,0.0000,-5220.8,-6268.9,-689.73,-1652.4,-817.09,-14556.,-84.792,-18277.,-5895.5,-3773.4,-2021.8,73.980,1641.6,1544.4,775.99,233.95,1579.9,1686.6,0.0000,5762.4,4449.7,4252.8,3658.0,0.0000,-223.71,-69.946,-47.977,-30.190,-30.751,-587.69,0.0000,-1038.1,-1490.5,-731.95,-1134.2
2018.000000000,61.594,1377.1,1394.8,740.86,197.27,1498.4,966.39,2.4132,4732.0,2763.1,3378.7,2119.4,0.0000,-5219.0,-6268.7,-688.32,-1651.9,-812.74,-14554.,-84.771,-18274.,-5895.2,-3773.0,-2021.4,45.543,1622.4,1479.4,774.72,222.31,1572.3,1686.6,0.0000,5757.7,4449.7,4252.8,3658.0,0.0000,-225.50,-68.862,-48.131,-30.362,-30.563,-587.69,0.0000,-1038.1,-1490.5,-731.93,-1134.1
2019.000000000,62.109,1387.9,1404.9,740.84,199.03,1494.1,966.39,2.4134,4728.1,2763.1,3378.7,2119.5,0.0000,-5217.6,-6268.8,-686.95,-1651.5,-808.45,-14553.,-84.749,-18272.,-5894.9,-3772.7,-2021.0,45.654,1626.4,1483.0,772.11,222.78,1564.3,1686.6,0.0000,5752.8,4449.7,4252.8,3658.0,0.0000,-226.00,-69.023,-48.101,-30.436,-30.369,-587.69,0.0000,-1038.0,-1490.4,-731.91,-1134.0
2020.000000000,62.526,1394.8,1411.9,740.62,200.09,1489.3,966.39,2.4137,4724.1,2763.1,3378.8,2119.6,0.0000,-5216.5,-6269.0,-685.64,-1651.0,-804.17,-14551.,-84.727,-18270.,-5894.6,-3772.3,-2020.7,45.662,1626.7,1483.3,768.99,222.76,1556.1,1686.6,0.0000,5747.8,4449.7,4252.8,3658.0,0.0000,-226.00,-69.030,-48.001,-30.442,-30.172,-587.69,0.0000,-1038.0,-1490.4,-731.88,-1133.9
2021.000000000,62.747,1398.2,1415.9,740.23,200.95,1484.0,966.39,2.4139,4720.0,2762.9,3378.8,2119.6,0.0000,-5215.5,-6269.1,-684.36,-1650.6,-799.87,-14549.,-84.705,-18268.,-5894.3,-3772.0,-2020.3,45.620,1625.2,1481.9,765.64,222.51,1547.8,1686.6,0.0000,5742.8,4449.7,4252.8,3658.0,0.0000,-225.74,-68.960,-47.867,-30.413,-29.976,-587.69,0.0000,-1038.0,-1490.3,-731.86,-1133.8
2022.000000000,62.952,1399.4,1417.5,739.15,201.35,1478.0,966.39,2.4141,4715.9,2762.9,3378.8,2119.7,0.0000,-5214.3,-6269.1,-683.13,-1650.1,-795.54,-14547.,-84.682,-18266.,-5894.0,-3771.6,-2019.9,45.545,1622.5,1479.5,762.13,222.10,1539.6,1686.6,0.0000,5737.8,4449.7,4252.8,3658.0,0.0000,-225.32,-68.840,-47.711,-30.363,-29.779,-587.69,0.0000,-1038.0,-1490.3,-731.83,-1133.8
2023.000000000,62.997,1399.3,1417.9,737.42,201.29,1471.6,966.39,2.4143,4711.6,2762.9,3378.7,2119.8,0.0000,-5213.1,-6269.0,-681.94,-1649.6,-791.18,-14546.,-84.660,-18263.,-5893.7,-3771.3,-2019.5,45.450,1619.1,1476.4,758.54,221.61,1531.3,1686.6,0.0000,5732.8,4449.7,4252.8,3658.0,0.0000,-224.81,-68.690,-47.543,-30.300,-29.583,-587.69,0.0000,-1038.0,-1490.2,-731.81,-1133.7
2024.000000000,62.953,1398.3,1417.4,735.40,201.02,1465.0,966.38,2.4145,4707.7,2763.0,3378.7,2119.9,0.0000,-5211.7,-6268.7,-680.79,-1649.1,-786.79,-14544.,-84.637,-18261.,-5893.3,-3770.9,-2019.2,45.344,1615.4,1473.0,754.93,221.06,1523.1,1686.6,0.0000,5727.8,4449.7,4252.8,3658.0,0.0000,-224.24,-68.522,-47.367,-30.230,-29.389,-587.69,0.0000,-1037.9,-1490.2,-731.79,-1133.6
2025.000000000,62.947,1397.1,1416.4,733.08,200.62,1457.8,966.36,2.4217,4704.3,2763.0,3378.7,2120.0,0.0000,-5210.1,-6268.3,-679.69,-1648.5,-782.38,-14542.,-84.614,-18259.,-5893.0,-3770.6,-2018.8,45.227,1611.2,1469.1,751.25,220.46,1514.9,1686.6,0.0000,5722.8,4449.7,4252.8,3658.0,0.0000,-223.62,-68.336,-47.184,-30.151,-29.194,-587.69,0.0000,-1037.9,-1490.1,-731.76,-1133.5
2026.000000000,62.867,1395.4,1415.1,730.58,200.16,1450.9,966.36,2.4437,4700.9,2763.1,3378.8,2120.1,0.0000,-5208.4,-6267.9,-678.64,-1647.9,-777.95,-14540.,-84.592,-18257.,-5892.7,-3770.2,-2018.4,45.100,1606.7,1465.0,747.51,219.81,1506.6,1686.6,0.0000,5717.8,4449.7,4252.8,3658.0,0.0000,-222.94,-68.135,-46.994,-30.067,-28.998,-587.69,0.0000,-1037.9,-1490.1,-731.74,-1133.4
2027.000000000,62.759,1393.0,1413.0,727.80,199.65,1444.3,966.36,2.4439,4698.3,2763.1,3378.8,2120.2,0.0000,-5206.6,-6267.3,-677.65,-1647.4,-773.50,-14539.,-84.569,-18255.,-5892.4,-3769.9,-2018.0,44.968,1602.0,1460.7,743.77,219.14,1498.4,1686.6,0.0000,5712.8,4449.7,4252.8,3658.0,0.0000,-222.24,-67.926,-46.800,-29.979,-28.803,-587.69,0.0000,-1037.9,-1490.0,-731.72,-1133.3
2028.000000000,62.640,1390.4,1410.3,724.99,199.11,1438.3,966.36,2.4442,4695.8,2763.2,3378.8,2120.3,0.0000,-5204.6,-6266.6,-676.74,-1646.8,-769.03,-14537.,-84.546,-18252.,-5892.1,-3769.5,-2017.6,44.835,1597.2,1456.4,740.05,218.47,1490.2,1686.6,0.0000,5707.9,4449.7,4252.8,3658.0,0.0000,-221.54,-67.714,-46.607,-29.890,-28.611,-587.69,0.0000,-1037.8,-1490.0,-731.69,-1133.2
2029.000000000,62.502,1387.3,1407.2,722.09,198.54,1432.9,966.36,2.4444,4693.3,2763.2,3378.8,2120.4,0.0000,-5202.5,-6265.9,-675.90,-1646.1,-764.53,-14535.,-84.523,-18250.,-5891.8,-3769.2,-2017.3,44.702,1592.5,1452.1,736.38,217.80,1482.2,1686.6,0.0000,5703.0,4449.7,4252.8,3658.0,0.0000,-220.83,-67.502,-46.416,-29.801,-28.420,-587.69,0.0000,-1037.8,-1489.9,-731.67,-1133.1
2030.000000000,62.371,1384.4,1403.8,718.99,197.97,1427.3,966.36,2.4446,4690.5,2763.2,3378.8,2120.5,0.0000,-5200.2,-6265.0,-675.18,-1645.5,-760.00,-14533.,-84.501,-18248.,-5891.5,-3768.8,-2016.9,44.566,1587.6,1447.7,732.69,217.11,1474.1,1686.6,0.0000,5698.2,4449.7,4252.8,3658.0,0.0000,-220.11,-67.283,-46.222,-29.711,-28.230,-587.69,0.0000,-1037.8,-1489.9,-731.64,-1133.0
2031.000000000,62.238,1381.3,1400.4,715.78,197.38,1421.7,966.36,2.4448,4687.2,2763.3,3378.9,2120.6,0.0000,-5197.7,-6264.2,-674.56,-1644.9,-755.44,-14532.,-84.478,-18246.,-5891.2,-3768.5,-2016.5,44.426,1582.7,1443.1,728.98,216.40,1466.1,1686.6,0.0000,5693.3,4449.7,4252.8,3658.0,0.0000,-219.37,-67.060,-46.025,-29.617,-28.039,-587.69,0.0000,-1037.8,-1489.8,-731.62,-1132.9
2032.000000000,62.102,1378.1,1397.2,712.56,196.78,1415.2,966.36,2.4450,4683.5,2763.3,3378.9,2120.7,0.0000,-5195.1,-6263.3,-674.07,-1644.3,-750.86,-14530.,-84.455,-18244.,-5890.9,-3768.1,-2016.1,44.288,1577.7,1438.6,725.30,215.70,1458.1,1686.6,0.0000,5688.5,4449.7,4252.8,3658.0,0.0000,-218.63,-66.838,-45.831,-29.525,-27.850,-587.69,0.0000,-1037.7,-1489.8,-731.60,-1132.8
2033.000000000,62.109,1374.7,1394.0,709.47,196.17,1408.4,966.36,2.4452,4679.5,2763.4,3378.9,2120.8,0.0000,-5192.4,-6262.3,-673.70,-1643.7,-746.24,-14528.,-84.433,-18242.,-5890.5,-3767.8,-2015.8,44.159,1573.1,1434.4,721.80,215.05,1450.4,1686.6,0.0000,5683.8,4449.7,4252.8,3658.0,0.0000,-217.94,-66.630,-45.646,-29.439,-27.667,-587.69,0.0000,-1037.7,-1489.7,-731.57,-1132.8
2034.000000000,62.014,1371.2,1390.7,706.30,195.59,1401.2,966.36,2.4455,4675.3,2763.4,3379.0,2120.9,0.0000,-5189.6,-6261.3,-673.45,-1643.0,-741.58,-14526.,-84.410,-18239.,-5890.2,-3767.4,-2015.4,44.036,1568.8,1430.4,718.39,214.43,1443.0,1686.6,0.0000,5679.3,4449.7,4252.8,3658.0,0.0000,-217.28,-66.431,-45.468,-29.357,-27.489,-587.69,0.0000,-1037.7,-1489.7,-731.55,-1132.7
2035.000000000,61.883,1367.8,1387.5,703.09,195.03,1393.7,966.36,2.4457,4671.0,2763.5,3379.0,2121.0,0.0000,-5186.8,-6260.2,-673.29,-1642.4,-736.90,-14525.,-84.388,-18237.,-5889.9,-3767.1,-2015.0,43.915,1564.5,1426.5,715.03,213.82,1435.6,1686.6,0.0000,5674.9,4449.7,4252.8,3658.0,0.0000,-216.63,-66.235,-45.292,-29.277,-27.313,-587.69,0.0000,-1037.7,-1489.6,-731.53,-1132.6
2036.000000000,61.754,1364.5,1384.4,699.83,194.47,1386.3,966.34,2.4483,4666.5,2763.5,3379.0,2121.1,0.0000,-5183.9,-6259.2,-673.18,-1641.7,-732.18,-14523.,-84.365,-18235.,-5889.6,-3766.7,-2014.6,43.792,1560.1,1422.5,711.65,213.19,1428.2,1686.6,0.0000,5670.4,4449.7,4252.8,3658.0,0.0000,-215.96,-66.034,-45.111,-29.194,-27.136,-587.69,0.0000,-1037.7,-1489.6,-731.50,-1132.5
2037.000000000,61.617,1361.1,1381.0,696.53,193.92,1378.9,966.32,2.4604,4662.1,2763.6,3379.0,2121.2,0.0000,-5181.0,-6258.0,-673.07,-1641.0,-727.43,-14521.,-84.342,-18233.,-5889.3,-3766.4,-2014.3,43.661,1555.4,1418.3,708.18,212.53,1420.7,1686.6,0.0000,5665.8,4449.7,4252.8,3658.0,0.0000,-215.26,-65.822,-44.920,-29.107,-26.956,-587.69,0.0000,-1037.6,-1489.5,-731.48,-1132.4
2038.000000000,61.490,1362.1,1380.9,693.29,193.88,1372.0,966.32,2.4606,4657.5,2763.6,3379.0,2121.3,0.0000,-5178.3,-6257.0,-672.99,-1640.4,-722.68,-14519.,-84.322,-18231.,-5889.0,-3766.0,-2013.9,63.480,1622.3,1477.1,727.92,222.69,1452.9,1686.6,9.1737,5685.4,4451.8,4256.3,3660.8,0.0000,-221.57,-68.112,-46.088,-29.987,-27.506,-587.69,-0.41886,-1037.6,-1489.5,-731.47,-1132.3
2039.000000000,61.623,1374.6,1391.0,690.67,196.27,1366.7,966.32,2.4608,4653.4,2763.7,3379.1,2121.3,0.0000,-5176.5,-6256.7,-672.96,-1639.9,-717.97,-14518.,-84.302,-18229.,-5888.7,-3765.7,-2013.5,45.592,1624.2,1481.0,729.16,221.74,1449.9,1686.6,0.0000,5684.2,4450.2,4254.5,3659.2,0.0000,-224.69,-68.715,-46.501,-30.395,-27.459,-587.69,0.0000,-1037.6,-1489.4,-731.44,-1132.2
2040.000000000,62.315,1388.9,1403.2,689.34,197.82,1362.4,966.31,2.4611,4650.0,2763.7,3379.1,2121.4,0.0000,-5175.4,-6256.8,-672.95,-1639.5,-713.28,-14516.,-84.282,-18227.,-5888.4,-3765.3,-2013.1,45.714,1628.5,1484.9,726.23,222.26,1443.0,1686.6,0.0000,5679.4,4449.9,4253.4,3658.5,0.0000,-225.25,-68.894,-46.493,-30.476,-27.303,-587.69,0.0000,-1037.6,-1489.4,-731.41,-1132.1
2041.000000000,62.619,1398.0,1412.3,689.17,198.39,1358.8,966.29,2.4613,4646.5,2763.4,3379.1,2121.5,0.0000,-5174.7,-6257.2,-672.94,-1639.1,-708.64,-14514.,-84.260,-18224.,-5888.1,-3765.0,-2012.8,45.724,1628.9,1485.3,723.26,222.26,1436.1,1686.6,0.0000,5675.0,4449.7,4253.0,3658.1,0.0000,-225.26,-68.906,-46.406,-30.483,-27.140,-587.69,0.0000,-1037.5,-1489.4,-731.38,-1132.0
2042.000000000,62.747,1402.3,1416.7,690.18,199.74,1356.0,966.30,2.4559,4643.2,2763.5,3379.1,2121.6,0.0000,-5174.0,-6257.6,-672.92,-1638.7,-704.05,-14512.,-84.239,-18222.,-5887.8,-3764.6,-2012.4,45.682,1627.4,1483.9,720.33,222.02,1429.3,1686.6,0.0000,5670.7,4449.7,4252.8,3658.0,0.0000,-225.02,-68.838,-46.282,-30.454,-26.976,-587.69,0.0000,-1037.5,-1489.3,-731.36,-1131.9
2043.000000000,63.136,1403.7,1418.2,690.30,200.61,1352.5,966.30,2.4609,4640.2,2763.5,3379.2,2121.7,0.0000,-5173.4,-6257.8,-672.90,-1638.3,-699.53,-14511.,-84.217,-18220.,-5887.4,-3764.3,-2012.0,45.609,1624.8,1481.5,717.37,221.63,1422.5,1686.6,0.0000,5666.6,4449.7,4252.8,3658.0,0.0000,-224.62,-68.723,-46.138,-30.406,-26.813,-587.69,0.0000,-1037.5,-1489.3,-731.34,-1131.8
2044.000000000,63.263,1403.6,1419.1,689.14,200.67,1348.1,966.30,2.4715,4636.8,2763.6,3379.2,2121.8,0.0000,-5172.6,-6257.8,-672.86,-1637.8,-694.98,-14509.,-84.194,-18218.,-5887.1,-3763.9,-2011.7,45.523,1621.7,1478.7,714.42,221.19,1415.9,1686.6,0.0000,5662.5,4449.7,4252.8,3658.0,0.0000,-224.16,-68.588,-45.986,-30.348,-26.652,-587.69,0.0000,-1037.5,-1489.2,-731.31,-1131.8
2045.000000000,63.238,1402.7,1418.4,688.02,200.42,1343.2,966.30,2.4718,4633.3,2763.6,3379.2,2121.8,0.0000,-5171.6,-6257.7,-672.82,-1637.3,-690.38,-14507.,-84.172,-18216.,-5886.8,-3763.6,-2011.3,45.421,1618.1,1475.4,711.40,220.67,1409.2,1686.6,0.0000,5658.5,4449.7,4252.8,3658.0,0.0000,-223.62,-68.429,-45.824,-30.281,-26.490,-587.69,0.0000,-1037.4,-1489.2,-731.29,-1131.7
2046.000000000,63.174,1401.1,1417.0,687.25,200.06,1337.8,966.30,2.4720,4629.8,2763.7,3379.2,2121.9,0.0000,-5170.5,-6257.5,-672.77,-1636.8,-685.75,-14505.,-84.150,-18214.,-5886.5,-3763.2,-2010.9,45.308,1614.1,1471.8,708.31,220.10,1402.4,1686.6,0.0000,5654.4,4449.7,4252.8,3658.0,0.0000,-223.02,-68.252,-45.653,-30.205,-26.328,-587.69,0.0000,-1037.4,-1489.1,-731.27,-1131.6
2047.000000000,63.085,1398.9,1416.0,685.61,199.62,1332.3,966.30,2.4722,4626.3,2763.7,3379.2,2122.0,0.0000,-5169.2,-6257.2,-672.72,-1636.3,-681.10,-14504.,-84.127,-18212.,-5886.2,-3762.9,-2010.5,45.187,1609.8,1467.8,705.17,219.49,1395.6,1686.6,0.0000,5650.3,4449.7,4252.8,3658.0,0.0000,-222.39,-68.063,-45.477,-30.125,-26.165,-587.69,0.0000,-1037.4,-1489.1,-731.24,-1131.5
2048.000000000,62.981,1396.3,1414.8,683.66,199.13,1326.9,966.30,2.4725,4623.0,2763.7,3379.3,2122.0,0.0000,-5167.9,-6256.8,-672.65,-1635.8,-676.43,-14502.,-84.105,-18210.,-5885.9,-3762.5,-2010.2,45.072,1605.7,1464.1,702.12,218.91,1389.0,1686.6,0.0000,5646.3,4449.7,4252.8,3658.0,0.0000,-221.79,-67.882,-45.308,-30.048,-26.006,-587.69,0.0000,-1037.4,-1489.0,-731.22,-1131.4
2049.000000000,62.870,1396.9,1415.5,681.19,198.93,1321.1,966.30,2.4727,4620.3,2763.8,3379.3,2122.1,0.0000,-5166.6,-6256.4,-672.60,-1635.2,-671.76,-14500.,-84.083,-18207.,-5885.6,-3762.2,-2009.8,98.488,1676.1,1504.1,708.81,225.20,1391.3,1686.6,0.0000,5647.0,4449.7,4252.8,3658.0,0.0000,-224.63,-69.192,-45.680,-30.452,-25.998,-587.69,0.0000,-1037.4,-1489.0,-731.19,-1131.3
2050.000000000,63.003,1402.7,1420.2,679.57,199.93,1315.2,966.30,2.4729,4617.0,2763.8,3379.4,2122.2,0.0000,-5165.7,-6256.2,-672.57,-1634.7,-667.10,-14498.,-84.063,-18205.,-5885.3,-3761.8,-2009.4,45.993,1669.0,1505.6,711.48,227.96,1391.0,1686.6,16.748,5649.4,4451.6,4255.2,3660.1,0.0000,-226.29,-69.505,-45.897,-30.691,-25.968,-587.69,-0.76468,-1037.4,-1488.9,-731.18,-1131.2
2051.000000000,63.378,1410.2,1426.8,678.23,200.77,1310.4,966.30,2.4732,4614.9,2763.9,3379.4,2122.3,0.0000,-5165.2,-6256.3,-672.56,-1634.3,-662.44,-14497.,-84.042,-18203.,-5885.0,-3761.5,-2009.0,103.24,1693.6,1547.2,718.25,242.55,1400.3,1686.6,38.311,5655.8,4457.8,4263.5,3668.5,0.0000,-227.89,-70.654,-46.130,-30.991,-26.021,-587.69,-1.7493,-1037.4,-1488.9,-731.20,-1131.2
2052.000000000,63.569,1418.3,1434.1,677.44,201.60,1306.6,966.30,2.4734,4613.4,2763.9,3379.4,2122.4,0.0000,-5165.0,-6256.7,-672.56,-1633.9,-657.79,-14495.,-84.022,-18201.,-5884.7,-3761.1,-2008.7,46.563,1658.8,1512.5,708.99,225.87,1390.0,1686.6,0.0000,5646.6,4449.7,4252.8,3658.0,0.0000,-228.99,-70.109,-46.243,-31.042,-25.905,-587.69,0.0000,-1037.3,-1488.8,-731.12,-1131.0
2053.000000000,63.846,1425.6,1440.6,676.95,202.71,1304.4,966.30,2.4736,4612.1,2764.0,3379.4,2122.4,0.0000,-5165.0,-6257.2,-672.57,-1633.6,-653.18,-14493.,-84.001,-18199.,-5884.4,-3760.8,-2008.3,46.585,1659.6,1513.3,707.02,225.94,1384.6,1686.6,0.0000,5643.3,4449.7,4252.8,3658.0,0.0000,-229.07,-70.142,-46.178,-31.057,-25.771,-587.69,0.0000,-1037.3,-1488.8,-731.10,-1131.0
2054.000000000,64.147,1429.5,1444.9,676.38,203.36,1302.0,966.30,2.4739,4610.4,2763.8,3379.4,2122.5,0.0000,-5165.0,-6257.7,-672.57,-1633.2,-648.59,-14491.,-83.980,-18197.,-5884.1,-3760.4,-2007.9,46.544,1658.1,1511.9,704.63,225.71,1378.9,1686.6,0.0000,5639.9,4449.7,4252.8,3658.0,0.0000,-228.84,-70.078,-46.068,-31.029,-25.630,-587.69,0.0000,-1037.2,-1488.7,-731.08,-1130.9
2055.000000000,64.265,1430.5,1446.9,675.54,203.69,1300.2,966.30,2.4377,4608.6,2763.7,3379.4,2122.6,0.0000,-5164.9,-6258.1,-672.56,-1632.9,-644.02,-14490.,-83.958,-18195.,-5883.8,-3760.1,-2007.6,46.467,1655.4,1509.4,702.03,225.31,1373.0,1686.6,0.0000,5636.3,4449.7,4252.8,3658.0,0.0000,-228.43,-69.961,-45.932,-30.978,-25.486,-587.69,0.0000,-1037.2,-1488.7,-731.05,-1130.8
2056.000000000,64.325,1430.3,1446.9,674.24,203.74,1297.3,966.30,2.2026,4606.3,2763.8,3379.5,2122.7,0.0000,-5164.7,-6258.4,-672.54,-1632.5,-639.47,-14488.,-83.936,-18193.,-5883.5,-3759.7,-2007.2,46.368,1651.8,1506.2,699.29,224.81,1367.0,1686.6,0.0000,5632.7,4449.7,4252.8,3658.0,0.0000,-227.92,-69.809,-45.780,-30.912,-25.340,-587.69,0.0000,-1037.2,-1488.6,-731.03,-1130.7
2057.000000000,64.053,1429.0,1446.2,672.81,203.51,1292.9,966.30,2.2078,4604.1,2763.8,3379.5,2122.8,0.0000,-5164.4,-6258.5,-672.52,-1632.1,-634.90,-14486.,-83.914,-18191.,-5883.2,-3759.4,-2006.8,46.255,1647.8,1502.5,696.48,224.24,1361.0,1686.6,0.0000,5629.0,4449.7,4252.8,3658.0,0.0000,-227.33,-69.637,-45.619,-30.837,-25.194,-587.69,0.0000,-1037.2,-1488.6,-731.01,-1130.6
2058.000000000,63.982,1427.3,1445.9,671.40,203.16,1288.4,966.31,2.2080,4601.3,2763.9,3379.5,2122.8,0.0000,-5163.9,-6258.6,-672.49,-1631.6,-630.32,-14484.,-83.892,-18189.,-5882.9,-3759.0,-2006.4,46.226,1646.8,1501.6,694.98,224.08,1357.4,1686.6,0.0000,5626.9,4449.7,4252.8,3658.0,0.0000,-227.16,-69.589,-45.542,-30.817,-25.097,-587.69,0.0000,-1037.1,-1488.5,-730.98,-1130.5
2059.000000000,63.904,1426.1,1445.1,669.74,202.91,1283.7,966.31,2.2082,4598.4,2763.9,3379.5,2122.9,0.0000,-5163.4,-6258.5,-672.45,-1631.2,-625.74,-14483.,-83.871,-18187.,-5882.5,-3758.7,-2006.1,46.192,1645.6,1504.1,694.76,236.82,1360.7,1686.6,0.0000,5626.8,4449.7,4252.8,3658.0,0.0000,-226.96,-69.612,-45.501,-30.874,-25.082,-587.69,0.0000,-1037.1,-1488.5,-730.96,-1130.4
2060.000000000,63.899,1425.6,1444.3,668.02,202.61,1279.0,966.31,2.2084,4595.6,2764.0,3379.5,2123.0,0.0000,-5162.8,-6258.4,-672.41,-1630.7,-621.16,-14481.,-83.849,-18185.,-5882.2,-3758.3,-2005.7,46.065,1641.0,1496.4,691.99,223.29,1351.5,1686.6,0.0000,5623.3,4449.7,4252.8,3658.0,0.0000,-226.31,-69.338,-45.335,-30.710,-24.927,-587.69,0.0000,-1037.1,-1488.5,-730.93,-1130.3
2061.000000000,63.915,1423.7,1442.6,666.51,202.14,1274.3,966.31,2.2086,4592.7,2764.0,3379.6,2123.1,0.0000,-5162.0,-6258.3,-672.37,-1630.2,-616.59,-14479.,-83.828,-18183.,-5881.9,-3758.0,-2005.3,45.935,1636.4,1492.1,689.18,222.64,1345.6,1686.6,0.0000,5619.8,4449.7,4252.8,3658.0,0.0000,-225.64,-69.136,-45.165,-30.623,-24.786,-587.69,0.0000,-1037.1,-1488.4,-730.91,-1130.2
2062.000000000,63.802,1421.0,1440.0,664.95,201.70,1269.7,966.31,2.2088,4589.8,2764.1,3379.6,2123.2,0.0000,-5161.0,-6258.0,-672.32,-1629.7,-612.03,-14478.,-83.806,-18180.,-5881.6,-3757.6,-2005.0,45.802,1631.7,1487.8,686.35,221.99,1339.8,1686.6,0.0000,5616.2,4449.7,4252.8,3658.0,0.0000,-224.95,-68.929,-44.993,-30.535,-24.645,-587.69,0.0000,-1037.0,-1488.4,-730.89,-1130.1
2063.000000000,63.703,1418.1,1436.6,663.35,201.28,1265.2,966.31,2.2090,4587.2,2764.1,3379.6,2123.3,0.0000,-5159.8,-6257.6,-672.27,-1629.2,-607.49,-14476.,-83.784,-18178.,-5881.3,-3757.3,-2004.6,45.669,1626.9,1483.5,683.54,221.33,1334.0,1686.6,0.0000,5612.7,4449.7,4252.8,3658.0,0.0000,-224.27,-68.722,-44.822,-30.446,-24.504,-587.69,0.0000,-1037.0,-1488.3,-730.86,-1130.1
2064.000000000,63.591,1415.1,1433.2,661.54,200.74,1260.9,966.31,2.2092,4584.9,2764.2,3379.7,2123.3,0.0000,-5158.5,-6257.1,-672.21,-1628.7,-602.96,-14474.,-83.762,-18176.,-5881.0,-3756.9,-2004.2,45.538,1622.3,1479.2,680.75,220.68,1328.2,1686.6,0.0000,5609.2,4449.7,4252.8,3658.0,0.0000,-223.58,-68.515,-44.652,-30.358,-24.365,-587.69,0.0000,-1037.0,-1488.3,-730.84,-1130.0
2065.000000000,63.398,1411.8,1429.9,659.50,200.10,1256.7,966.31,2.2094,4582.9,2764.2,3379.7,2123.3,0.0000,-5157.0,-6256.5,-672.16,-1628.2,-598.42,-14472.,-83.740,-18174.,-5880.7,-3756.6,-2003.9,45.406,1617.6,1475.0,677.97,220.03,1322.5,1686.6,0.0000,5605.8,4449.7,4252.8,3658.0,0.0000,-222.90,-68.309,-44.483,-30.271,-24.227,-587.69,0.0000,-1037.0,-1488.2,-730.82,-1129.9
2066.000000000,63.172,1408.5,1426.2,657.18,199.54,1252.7,966.31,2.2096,4580.8,2764.3,3379.7,2123.4,0.0000,-5155.3,-6255.8,-672.09,-1627.6,-593.88,-14471.,-83.718,-18172.,-5880.4,-3756.2,-2003.5,45.275,1612.9,1470.7,675.21,219.38,1316.8,1686.6,0.0000,5602.3,4449.7,4252.8,3658.0,0.0000,-222.22,-68.102,-44.315,-30.183,-24.090,-587.69,0.0000,-1037.0,-1488.2,-730.79,-1129.8
2067.000000000,62.980,1405.2,1422.7,655.13,198.98,1249.2,966.31,2.2098,4578.6,2764.3,3379.7,2123.5,0.0000,-5153.5,-6255.1,-672.03,-1627.1,-589.32,-14469.,-83.696,-18170.,-5880.1,-3755.9,-2003.1,45.144,1608.2,1466.4,672.45,218.73,1311.1,1686.6,0.0000,5598.9,4449.7,4252.8,3658.0,0.0000,-221.53,-67.895,-44.147,-30.096,-23.953,-587.69,0.0000,-1036.9,-1488.1,-730.77,-1129.7
2068.000000000,62.844,1401.7,1419.7,652.59,198.42,1245.0,966.31,2.2100,4576.0,2764.4,3379.7,2123.6,0.0000,-5151.6,-6254.3,-671.96,-1626.5,-584.77,-14467.,-83.674,-18168.,-5879.8,-3755.5,-2002.7,45.014,1603.6,1462.2,669.72,218.09,1305.5,1686.6,0.0000,5595.5,4449.7,4252.8,3658.0,0.0000,-220.85,-67.689,-43.981,-30.010,-23.818,-587.69,0.0000,-1036.9,-1488.1,-730.75,-1129.6
2069.000000000,62.712,1398.1,1416.7,650.15,197.85,1240.6,966.31,2.2102,4573.2,2764.4,3379.8,2123.7,0.0000,-5149.6,-6253.5,-671.90,-1625.9,-580.21,-14465.,-83.652,-18166.,-5879.5,-3755.2,-2002.4,44.886,1599.1,1458.1,667.02,217.45,1299.9,1686.6,0.0000,5592.1,4449.7,4252.8,3658.0,0.0000,-220.18,-67.486,-43.816,-29.924,-23.684,-587.69,0.0000,-1036.9,-1488.0,-730.72,-1129.5
