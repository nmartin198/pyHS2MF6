time,RECHARGE,RECHARGE,RECHARGE,RECHARGE,RECHARGE,RECHARGE,RECHARGE,RECHARGE,RECHARGE,RECHARGE,RECHARGE,RECHARGE,DISCHARGE,DISCHARGE,DISCHARGE,DISCHARGE,DISCHARGE,DISCHARGE,DISCHARGE,DISCHARGE,DISCHARGE,DISCHARGE,DISCHARGE,DISCHARGE,INFILT,INFILT,INFILT,INFILT,INFILT,INFILT,INFILT,INFILT,INFILT,INFILT,INFILT,INFILT,REJINFILT,REJINFILT,REJINFILT,REJINFILT,REJINFILT,REJINFILT,REJINFILT,REJINFILT,REJINFILT,REJINFILT,REJINFILT,REJINFILT
1.000000000000,0.62700E+06,0.10864E+06,0.13610E+06,0.13377E+06,0.16464E+06,91843.,0.22563E+06,35976.,0.13025E+06,26687.,54288.,62806.,0.0000,-3978.9,-6953.1,-321.89,-2380.2,-3205.5,-13851.,-1665.8,-1701.0,-5218.8,-2523.9,-5724.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
2.000000000000,0.62628E+06,0.10611E+06,0.13453E+06,0.13353E+06,0.16316E+06,90843.,0.22345E+06,35496.,0.12959E+06,26172.,53186.,61947.,0.0000,-4127.5,-7191.5,-328.92,-2503.2,-3274.9,-14350.,-1669.1,-1805.7,-5395.6,-2605.8,-5881.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
3.000000000000,0.62598E+06,0.10378E+06,0.13226E+06,0.13325E+06,0.16073E+06,89533.,0.22154E+06,35040.,0.12871E+06,25528.,52319.,60999.,0.0000,-4235.6,-7317.7,-337.50,-2604.1,-3331.5,-14813.,-1672.8,-1898.9,-5503.0,-2647.0,-6006.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
4.000000000000,0.62610E+06,0.10172E+06,0.13008E+06,0.13268E+06,0.15825E+06,87810.,0.22009E+06,34619.,0.12735E+06,24901.,51372.,60165.,0.0000,-4381.1,-7407.3,-351.14,-2686.5,-3409.6,-15203.,-1679.1,-2012.0,-5587.7,-2669.1,-6112.8,18857.,8428.7,6456.6,6059.7,11747.,4048.0,14510.,4193.0,6410.0,1913.3,2749.8,3312.2,0.0000,-21.641,-20.477,-3.0528,-19.183,-15.892,-76.664,-59.097,-6.1055,-53.658,-6.3452,-72.165
5.000000000000,0.62455E+06,99475.,0.12807E+06,0.13130E+06,0.15607E+06,85361.,0.21792E+06,34073.,0.12553E+06,24213.,50526.,59352.,0.0000,-4496.2,-7481.3,-364.98,-2748.5,-3464.3,-15520.,-1683.3,-2097.4,-5642.5,-2689.0,-6196.7,9936.3,4441.3,3402.2,3193.1,6189.9,2133.0,7645.6,2209.4,3377.6,1008.2,1448.9,1745.3,0.0000,-11.589,-10.868,-1.6086,-10.190,-8.5434,-40.967,-31.146,-3.2172,-28.315,-3.3449,-38.042
6.000000000000,0.62318E+06,97347.,0.12641E+06,0.12981E+06,0.15449E+06,82908.,0.21556E+06,33539.,0.12369E+06,23650.,49657.,58695.,0.0000,-4555.0,-7527.3,-373.95,-2799.1,-3496.9,-15785.,-1685.7,-2134.9,-5670.1,-2705.8,-6256.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
7.000000000000,0.62215E+06,95522.,0.12462E+06,0.12846E+06,0.15361E+06,80635.,0.21349E+06,32945.,0.12177E+06,23050.,48851.,58042.,0.0000,-4626.0,-7567.1,-382.14,-2844.0,-3557.5,-16009.,-1688.0,-2179.6,-5691.7,-2722.5,-6306.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
8.000000000000,0.62122E+06,93281.,0.12273E+06,0.12702E+06,0.15237E+06,77962.,0.21086E+06,32518.,0.11903E+06,22381.,48219.,57442.,0.0000,-4693.7,-7605.7,-389.93,-2881.8,-3618.3,-16198.,-1690.3,-2218.2,-5710.0,-2740.3,-6348.6,259.09,115.81,88.712,83.259,161.40,55.618,199.36,57.610,88.073,26.289,37.781,45.510,0.0000,-0.31265,-0.28822,-0.41944E-01,-0.27003,-0.23036,-1.1111,-0.81258,-0.83889E-01,-0.74079,-0.88329E-01,-0.99302
9.000000000000,0.62033E+06,91160.,0.12106E+06,0.12571E+06,0.15129E+06,75478.,0.20858E+06,32123.,0.11637E+06,21744.,47491.,56799.,0.0000,-4810.1,-7674.3,-401.75,-2912.8,-3718.5,-16403.,-1707.6,-2287.4,-5739.4,-2758.9,-6396.8,0.11223E+06,50164.,38427.,36065.,69914.,24092.,86357.,24955.,38150.,11387.,16366.,19713.,0.0000,-137.00,-125.48,-18.169,-117.71,-100.94,-485.86,-352.10,-36.338,-321.19,-38.428,-430.30
10.00000000000,0.61890E+06,88444.,0.11924E+06,0.12432E+06,0.14920E+06,73274.,0.20611E+06,31572.,0.11321E+06,21038.,46522.,55913.,0.0000,-4898.0,-7738.1,-413.25,-2943.3,-3793.9,-16627.,-1723.6,-2335.4,-5761.2,-2774.1,-6437.1,0.13078E+06,58456.,44779.,42026.,81470.,28074.,0.10063E+06,29080.,44456.,13270.,19071.,22972.,0.0000,-161.38,-146.92,-21.172,-137.93,-118.84,-571.29,-410.48,-42.344,-374.41,-44.962,-501.60
11.00000000000,0.61686E+06,86515.,0.11667E+06,0.12314E+06,0.14766E+06,71087.,0.20263E+06,31050.,0.11086E+06,20301.,45748.,54956.,0.0000,-4925.2,-7767.3,-419.51,-2974.1,-3813.8,-16816.,-1718.2,-2341.5,-5769.5,-2786.3,-6460.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
12.00000000000,0.61499E+06,85308.,0.11460E+06,0.12187E+06,0.14525E+06,69339.,0.19929E+06,30368.,0.10813E+06,19487.,44771.,53923.,0.0000,-4974.1,-7798.2,-424.81,-3005.5,-3850.1,-16963.,-1714.2,-2358.5,-5781.5,-2802.0,-6481.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
13.00000000000,0.61375E+06,82205.,0.11232E+06,0.12044E+06,0.14075E+06,67661.,0.19688E+06,29837.,0.10535E+06,18746.,43839.,52915.,0.0000,-5021.0,-7824.5,-430.14,-3037.7,-3882.6,-17079.,-1711.7,-2371.9,-5790.6,-2817.4,-6498.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
14.00000000000,0.60970E+06,79795.,0.11028E+06,0.11901E+06,0.13848E+06,65462.,0.19427E+06,29395.,0.10269E+06,18110.,42930.,51978.,0.0000,-5062.1,-7846.8,-434.62,-3069.1,-3909.0,-17187.,-1710.4,-2381.6,-5795.3,-2831.5,-6510.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
15.00000000000,0.60552E+06,77932.,0.10718E+06,0.11692E+06,0.13715E+06,64201.,0.19093E+06,28775.,0.10024E+06,17404.,42005.,51087.,0.0000,-5099.7,-7870.4,-438.55,-3098.4,-3930.2,-17291.,-1709.9,-2389.1,-5792.5,-2844.8,-6521.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
16.00000000000,0.60352E+06,75553.,0.10404E+06,0.11504E+06,0.13136E+06,62498.,0.18872E+06,28325.,97968.,16627.,41272.,50316.,0.0000,-5135.5,-7891.2,-442.35,-3120.7,-3948.8,-17377.,-1710.1,-2392.2,-5788.3,-2856.9,-6534.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
17.00000000000,0.59852E+06,73044.,0.10179E+06,0.11380E+06,0.12645E+06,60627.,0.18544E+06,27774.,94918.,16102.,40497.,49135.,0.0000,-5170.4,-7900.3,-446.12,-3140.9,-3964.7,-17451.,-1710.6,-2394.3,-5782.7,-2867.2,-6545.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
18.00000000000,0.59220E+06,70033.,99266.,0.11197E+06,0.12351E+06,59208.,0.18307E+06,27182.,91901.,15682.,39533.,47991.,0.0000,-5201.2,-7905.3,-449.84,-3160.4,-3976.4,-17517.,-1711.4,-2395.4,-5779.3,-2875.8,-6555.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
19.00000000000,0.58669E+06,67242.,96220.,0.10949E+06,0.12209E+06,58188.,0.18028E+06,26645.,90150.,15265.,38768.,47273.,0.0000,-5229.8,-7909.1,-453.48,-3179.7,-3985.8,-17579.,-1712.3,-2396.3,-5774.1,-2883.3,-6565.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
20.00000000000,0.58170E+06,63958.,93106.,0.10753E+06,0.11913E+06,56690.,0.17651E+06,26164.,88371.,14625.,38044.,46576.,0.0000,-5255.1,-7913.1,-456.89,-3195.0,-3993.3,-17628.,-1713.3,-2396.5,-5767.7,-2890.1,-6575.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
21.00000000000,0.57476E+06,61710.,90341.,0.10600E+06,0.11591E+06,55923.,0.17360E+06,25652.,86513.,14040.,37356.,45613.,0.0000,-5278.1,-7915.1,-459.54,-3206.6,-3997.0,-17667.,-1714.3,-2394.8,-5763.4,-2896.1,-6582.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
22.00000000000,0.56636E+06,58802.,86398.,0.10462E+06,0.11100E+06,54562.,0.17153E+06,24977.,83841.,13575.,36701.,44225.,0.0000,-5300.4,-7918.9,-461.89,-3217.6,-3997.9,-17700.,-1715.3,-2391.2,-5759.2,-2901.9,-6586.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
23.00000000000,0.56177E+06,56169.,83717.,0.10255E+06,0.10564E+06,53083.,0.16856E+06,24422.,81533.,13166.,35794.,42983.,0.0000,-5321.2,-7926.0,-464.15,-3227.9,-3997.9,-17724.,-1716.3,-2384.0,-5755.3,-2906.7,-6589.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
24.00000000000,0.55513E+06,53602.,81506.,0.10024E+06,0.10260E+06,51714.,0.16605E+06,23915.,79352.,12839.,35002.,42153.,0.0000,-5338.5,-7934.6,-466.37,-3238.7,-3995.8,-17743.,-1717.2,-2377.1,-5751.9,-2910.8,-6591.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
25.00000000000,0.54543E+06,50297.,79021.,98353.,96558.,50343.,0.16214E+06,23339.,77660.,12397.,33946.,41351.,0.0000,-5353.8,-7940.2,-468.55,-3250.0,-3992.4,-17757.,-1718.1,-2368.7,-5749.0,-2916.0,-6590.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
26.00000000000,0.53382E+06,46906.,76616.,96423.,93171.,49109.,0.15829E+06,22903.,75444.,12013.,32711.,40507.,0.0000,-5367.9,-7946.4,-470.41,-3261.2,-3988.2,-17768.,-1719.0,-2359.8,-5745.7,-2921.4,-6588.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
27.00000000000,0.52345E+06,45065.,74036.,94400.,91315.,48250.,0.15569E+06,22472.,73336.,11698.,31845.,39482.,0.0000,-5381.2,-7952.1,-472.00,-3272.3,-3982.2,-17778.,-1719.8,-2350.9,-5741.6,-2926.4,-6586.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
28.00000000000,0.51387E+06,42989.,70421.,91715.,87479.,47179.,0.15323E+06,22095.,71315.,11467.,31167.,38496.,0.0000,-5394.5,-7955.3,-473.50,-3283.3,-3974.6,-17785.,-1720.6,-2340.3,-5734.6,-2930.6,-6582.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
29.00000000000,0.50672E+06,41102.,67977.,89501.,83712.,45586.,0.14967E+06,21709.,69284.,11079.,30572.,37515.,0.0000,-5407.3,-7954.9,-474.96,-3293.9,-3966.5,-17781.,-1721.4,-2330.1,-5728.0,-2934.6,-6579.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
30.00000000000,0.49721E+06,39441.,66667.,86383.,80715.,44501.,0.14581E+06,21324.,67151.,10673.,29718.,36467.,0.0000,-5418.1,-7955.8,-476.40,-3299.9,-3958.4,-17763.,-1722.1,-2320.4,-5723.2,-2938.7,-6575.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
31.00000000000,0.47385E+06,38398.,65381.,84545.,75071.,43599.,0.14270E+06,21004.,64718.,10312.,28970.,35328.,0.0000,-5425.6,-7958.5,-477.81,-3305.0,-3950.7,-17740.,-1722.8,-2311.4,-5718.7,-2942.4,-6572.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
32.00000000000,0.45530E+06,36459.,63918.,81507.,69839.,42333.,0.13872E+06,20612.,62236.,9970.5,28198.,34034.,0.0000,-5432.2,-7962.7,-479.19,-3310.0,-3943.5,-17715.,-1723.4,-2302.8,-5714.4,-2945.6,-6568.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
33.00000000000,0.44015E+06,34458.,62291.,78604.,66921.,41455.,0.13387E+06,20142.,60062.,9769.2,27081.,32724.,0.0000,-5438.6,-7967.2,-480.55,-3315.1,-3936.1,-17690.,-1724.0,-2294.0,-5710.3,-2948.7,-6563.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
34.00000000000,0.42607E+06,32256.,60793.,77050.,65081.,40486.,0.13066E+06,19773.,57882.,9593.2,26145.,31923.,0.0000,-5444.0,-7971.5,-481.87,-3320.7,-3928.6,-17666.,-1724.5,-2284.9,-5706.3,-2952.1,-6559.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
35.00000000000,0.41863E+06,30985.,57606.,74964.,63466.,39759.,0.12819E+06,19466.,56348.,9469.8,25225.,31209.,0.0000,-5449.1,-7975.0,-483.15,-3326.2,-3921.2,-17639.,-1725.1,-2275.7,-5702.3,-2955.8,-6554.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
36.00000000000,0.41226E+06,28989.,55798.,72877.,61546.,38739.,0.12526E+06,19035.,54898.,9261.4,24514.,30348.,0.0000,-5453.2,-7978.3,-484.38,-3331.2,-3912.9,-17606.,-1725.6,-2266.1,-5698.0,-2959.5,-6549.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
37.00000000000,0.39749E+06,27764.,54510.,71862.,59163.,37721.,0.12045E+06,18761.,53310.,8906.9,23864.,29773.,0.0000,-5455.7,-7981.5,-485.51,-3336.4,-3903.9,-17573.,-1726.1,-2255.3,-5694.0,-2962.8,-6545.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
38.00000000000,0.38153E+06,26629.,53915.,70136.,57173.,37147.,0.11619E+06,18344.,52177.,8642.0,22859.,28870.,0.0000,-5458.1,-7983.7,-486.47,-3341.8,-3894.4,-17537.,-1726.6,-2243.8,-5690.0,-2965.5,-6541.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
39.00000000000,0.36716E+06,25850.,53251.,67671.,56225.,36204.,0.11363E+06,17900.,50400.,8344.3,21975.,27629.,0.0000,-5460.7,-7985.7,-487.00,-3347.1,-3884.5,-17501.,-1727.1,-2232.5,-5686.1,-2968.1,-6536.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
40.00000000000,0.34593E+06,25545.,51060.,65114.,55011.,35285.,0.11026E+06,17541.,48560.,8026.4,21399.,26600.,0.0000,-5463.6,-7988.0,-487.44,-3352.4,-3873.8,-17467.,-1727.5,-2221.4,-5681.3,-2970.3,-6530.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
41.00000000000,0.33451E+06,24640.,47952.,62652.,51941.,34370.,0.10634E+06,17194.,46748.,7751.3,20845.,25545.,0.0000,-5466.6,-7990.6,-487.85,-3358.0,-3862.7,-17432.,-1728.0,-2209.0,-5676.4,-2972.2,-6524.5,743.47,332.32,254.56,238.92,463.15,159.60,572.08,165.32,252.73,75.437,108.42,130.59,0.0000,-0.99778,-0.90526,-0.12036,-0.82141,-0.75521,-3.4829,-2.3502,-0.24072,-2.1403,-0.26969,-2.8600
42.00000000000,0.32245E+06,23640.,46791.,60589.,48608.,33344.,0.10315E+06,16805.,45919.,7549.7,20130.,24674.,0.0000,-5469.4,-7994.0,-488.24,-3363.8,-3851.1,-17399.,-1728.4,-2195.2,-5671.7,-2974.1,-6517.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
43.00000000000,0.31540E+06,23026.,46010.,58777.,47264.,32221.,99651.,16313.,44985.,7410.3,19404.,23973.,0.0000,-5472.0,-7998.6,-488.62,-3368.2,-3839.9,-17362.,-1728.7,-2180.1,-5667.3,-2976.2,-6510.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
44.00000000000,0.30825E+06,22447.,44280.,55970.,46358.,30922.,96425.,15920.,43028.,7311.6,18788.,23282.,0.0000,-5473.7,-8001.3,-489.00,-3372.6,-3829.4,-17321.,-1729.0,-2165.7,-5663.4,-2978.2,-6504.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
45.00000000000,0.29968E+06,21728.,41841.,54424.,44825.,29951.,93566.,15483.,42768.,7154.8,18186.,22619.,0.0000,-5472.9,-8001.5,-489.38,-3377.2,-3819.4,-17278.,-1729.3,-2152.0,-5660.0,-2980.2,-6497.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
46.00000000000,0.29268E+06,21128.,39472.,53399.,41148.,29414.,90876.,15213.,41384.,6953.5,17686.,21921.,0.0000,-5470.4,-7998.9,-489.77,-3381.8,-3809.9,-17227.,-1729.6,-2138.5,-5656.6,-2982.1,-6490.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
47.00000000000,0.27893E+06,20277.,38943.,52244.,38762.,28439.,87742.,14818.,40357.,6753.9,17159.,21337.,0.0000,-5467.2,-7995.7,-490.15,-3386.3,-3800.7,-17177.,-1729.8,-2125.3,-5652.8,-2984.0,-6483.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
48.00000000000,0.26751E+06,19602.,37987.,50478.,37752.,28103.,84169.,14261.,39173.,6595.5,16417.,20942.,0.0000,-5464.2,-7989.3,-490.53,-3390.7,-3791.1,-17130.,-1730.1,-2112.2,-5648.9,-2985.9,-6476.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
49.00000000000,0.25771E+06,18971.,37327.,48637.,36811.,27438.,81682.,13549.,37835.,6498.0,15784.,20481.,0.0000,-5461.0,-7982.9,-490.90,-3395.0,-3781.5,-17085.,-1730.3,-2099.4,-5645.6,-2987.8,-6469.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
50.00000000000,0.25317E+06,18168.,36754.,47000.,36274.,26860.,80081.,13236.,37050.,6270.7,15264.,19711.,0.0000,-5457.8,-7977.4,-491.22,-3399.1,-3771.5,-17043.,-1730.4,-2087.0,-5642.2,-2989.5,-6463.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
51.00000000000,0.25060E+06,17970.,34702.,45776.,35672.,26434.,77780.,12866.,36124.,6077.9,14832.,19248.,0.0000,-5454.4,-7970.4,-491.49,-3403.2,-3761.8,-17003.,-1730.6,-2075.1,-5638.9,-2991.0,-6457.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
52.00000000000,0.24539E+06,17683.,33308.,44658.,34907.,25662.,76196.,12580.,35919.,5934.2,14405.,18737.,0.0000,-5503.9,-7994.2,-496.10,-3407.5,-3797.4,-16967.,-1731.7,-2097.3,-5645.8,-2994.9,-6459.5,6393.2,2857.6,2189.0,2054.5,3982.7,1372.4,4919.4,1421.6,2173.2,648.69,932.28,1123.0,0.0000,-8.5959,-7.9341,-1.0350,-7.0911,-6.6213,-29.712,-20.240,-2.0700,-18.415,-2.3323,-24.601
53.00000000000,0.24076E+06,16908.,32913.,43341.,34100.,24648.,74615.,12196.,35034.,5781.4,14140.,18463.,0.0000,-5475.7,-7989.9,-495.90,-3411.5,-3766.8,-16931.,-1731.7,-2069.1,-5633.5,-2994.6,-6448.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
54.00000000000,0.23474E+06,16463.,32226.,42211.,32778.,23939.,72940.,11998.,34289.,5657.9,13918.,18197.,0.0000,-5467.5,-7981.9,-495.25,-3415.1,-3753.5,-16898.,-1731.7,-2054.7,-5627.9,-2995.5,-6441.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
55.00000000000,0.22866E+06,15958.,31846.,41505.,32175.,23217.,71062.,11747.,33612.,5398.3,13520.,17738.,0.0000,-5461.6,-7974.1,-494.74,-3416.6,-3742.7,-16861.,-1731.8,-2043.1,-5624.2,-2996.7,-6434.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
56.00000000000,0.22236E+06,15727.,31628.,39883.,30857.,22504.,68934.,11570.,32871.,5285.2,13145.,17149.,0.0000,-5509.3,-7997.4,-498.78,-3416.9,-3777.3,-16816.,-1732.8,-2065.8,-5632.9,-3000.7,-6437.1,6180.3,2762.5,2116.1,1986.1,3850.1,1326.7,4755.6,1374.2,2100.9,627.09,901.24,1085.6,0.0000,-8.3182,-7.7193,-1.0005,-6.8608,-6.4406,-28.624,-19.574,-2.0011,-17.803,-2.2577,-23.784
57.00000000000,0.21469E+06,15531.,31310.,39086.,29461.,21908.,67420.,11234.,31962.,5164.3,12802.,16583.,0.0000,-5479.2,-7992.2,-498.15,-3416.8,-3747.2,-16771.,-1732.7,-2038.5,-5621.8,-3000.5,-6426.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
58.00000000000,0.19966E+06,15272.,28561.,38404.,29018.,21126.,66421.,10995.,30630.,4995.4,12539.,16225.,0.0000,-5468.9,-7981.6,-497.08,-3416.7,-3734.4,-16727.,-1732.6,-2024.6,-5616.9,-3001.5,-6419.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
59.00000000000,0.19258E+06,14871.,28190.,37216.,28435.,20765.,64635.,10790.,29801.,4885.1,12246.,15624.,0.0000,-5460.9,-7971.7,-496.17,-3416.7,-3724.0,-16688.,-1732.6,-2012.6,-5613.5,-3002.7,-6413.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
60.00000000000,0.18857E+06,14584.,28052.,36134.,28033.,20118.,62802.,10411.,28854.,4698.5,11972.,14899.,0.0000,-5453.7,-7962.9,-495.46,-3416.8,-3714.7,-16647.,-1732.6,-2001.5,-5610.7,-3003.9,-6407.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
61.00000000000,0.18202E+06,14237.,27834.,34786.,27422.,19927.,60028.,10038.,28111.,4640.1,11710.,14473.,0.0000,-5447.1,-7955.0,-494.91,-3417.0,-3706.1,-16609.,-1732.6,-1991.3,-5608.2,-3005.1,-6402.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
62.00000000000,0.17735E+06,14023.,27411.,33808.,26799.,19566.,58548.,9564.6,27645.,4594.2,11421.,14062.,0.0000,-5440.9,-7948.1,-494.46,-3417.8,-3697.9,-16572.,-1732.7,-1981.8,-5606.0,-3006.4,-6396.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
63.00000000000,0.17249E+06,13683.,27264.,32981.,26510.,18917.,57144.,9318.7,27090.,4530.6,11116.,13958.,0.0000,-5434.9,-7942.0,-494.07,-3418.7,-3689.9,-16538.,-1732.8,-1972.9,-5603.9,-3007.7,-6390.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
64.00000000000,0.17014E+06,13427.,27019.,32298.,26225.,18453.,55865.,9121.9,26015.,4456.5,10711.,13749.,0.0000,-5428.9,-7936.9,-493.73,-3419.7,-3682.1,-16506.,-1732.9,-1963.9,-5601.8,-3009.1,-6384.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
65.00000000000,0.16751E+06,12980.,25182.,31291.,25803.,17893.,54961.,8855.5,25273.,4384.3,10466.,13413.,0.0000,-5422.9,-7932.3,-493.42,-3420.5,-3674.5,-16476.,-1733.0,-1954.9,-5599.7,-3010.4,-6378.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
66.00000000000,0.16606E+06,12505.,24028.,30367.,25486.,17624.,53832.,8637.4,25015.,4295.5,10179.,13140.,0.0000,-5416.9,-7928.0,-493.11,-3421.0,-3667.1,-16447.,-1733.1,-1945.9,-5597.7,-3011.7,-6373.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
67.00000000000,0.16510E+06,12193.,23675.,30043.,24994.,17188.,52784.,8453.2,24430.,4155.1,9949.1,12829.,0.0000,-5411.0,-7923.8,-492.81,-3421.6,-3660.1,-16418.,-1733.3,-1937.3,-5595.7,-3013.0,-6367.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
68.00000000000,0.16152E+06,11796.,23553.,29601.,24790.,16983.,51199.,8404.0,23842.,4067.3,9740.0,12596.,0.0000,-5405.1,-7919.8,-492.50,-3422.3,-3653.0,-16386.,-1733.4,-1928.8,-5593.7,-3014.2,-6362.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
69.00000000000,0.15671E+06,11639.,23111.,29407.,24196.,16768.,49665.,8309.0,23544.,3933.6,9624.6,12452.,0.0000,-5452.2,-7945.8,-496.58,-3423.4,-3686.5,-16355.,-1736.1,-1953.1,-5604.2,-3018.0,-6366.4,19330.,8640.1,6618.6,6211.8,12042.,4149.5,14874.,4298.2,6570.9,1961.3,2818.8,3395.3,0.0000,-25.851,-24.477,-3.1294,-21.429,-20.456,-88.547,-61.280,-6.2587,-55.681,-7.1416,-74.400
70.00000000000,0.15199E+06,11405.,22999.,29072.,23742.,16613.,47980.,8171.4,23260.,3778.5,9474.4,12276.,0.0000,-5421.8,-7945.0,-495.87,-3424.5,-3659.6,-16324.,-1735.6,-1928.3,-5594.7,-3017.4,-6356.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
71.00000000000,0.14755E+06,10996.,22912.,28610.,23241.,16427.,46661.,8019.9,22552.,3706.7,9226.5,12018.,0.0000,-5411.4,-7939.4,-494.75,-3425.5,-3649.0,-16294.,-1735.1,-1916.0,-5590.8,-3018.0,-6349.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
72.00000000000,0.14386E+06,10658.,22811.,27937.,23162.,15877.,45787.,7805.5,22224.,3657.3,9047.5,11808.,0.0000,-5403.4,-7933.0,-493.53,-3426.6,-3640.4,-16265.,-1734.9,-1905.7,-5588.0,-3018.8,-6343.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
73.00000000000,0.14219E+06,10595.,22421.,26892.,23005.,15578.,45338.,7708.1,21703.,3601.6,8923.7,11450.,0.0000,-5395.9,-7925.5,-492.44,-3427.7,-3632.4,-16237.,-1734.7,-1896.2,-5585.3,-3019.6,-6338.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
74.00000000000,0.14008E+06,10491.,22183.,26357.,22874.,15393.,44880.,7670.7,21128.,3511.1,8784.2,11265.,0.0000,-5388.4,-7918.6,-491.48,-3428.9,-3624.5,-16210.,-1734.5,-1887.0,-5582.6,-3020.5,-6332.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
75.00000000000,0.13764E+06,10342.,20341.,25978.,21492.,15102.,43967.,7591.1,20580.,3449.4,8691.4,11057.,0.0000,-5381.1,-7912.2,-490.62,-3430.1,-3616.7,-16184.,-1734.4,-1878.1,-5580.2,-3021.5,-6327.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
76.00000000000,0.13637E+06,9948.0,18543.,25304.,20911.,14919.,43149.,7450.5,20391.,3420.1,8558.5,10777.,0.0000,-5374.1,-7906.2,-489.83,-3431.4,-3609.1,-16158.,-1734.4,-1868.9,-5578.0,-3022.5,-6322.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
77.00000000000,0.13446E+06,9678.1,18127.,25125.,20855.,14670.,42583.,7358.9,20101.,3353.1,8417.3,10607.,0.0000,-5367.0,-7900.4,-489.09,-3432.8,-3601.8,-16134.,-1734.4,-1859.6,-5575.9,-3023.5,-6316.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
78.00000000000,0.13240E+06,9382.8,17891.,24687.,20634.,14164.,41886.,7250.0,19826.,3312.9,8260.8,10461.,0.0000,-5360.0,-7894.9,-488.38,-3434.1,-3594.7,-16110.,-1734.4,-1850.9,-5573.8,-3024.4,-6311.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
79.00000000000,0.13117E+06,9373.1,17737.,23945.,20235.,13796.,41135.,7086.6,19578.,3277.1,8114.0,10277.,0.0000,-5353.2,-7889.6,-487.70,-3435.6,-3588.0,-16087.,-1734.4,-1842.6,-5571.6,-3025.3,-6305.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
80.00000000000,0.13034E+06,9242.0,17480.,23687.,20072.,13678.,40534.,6931.4,19261.,3225.7,7976.0,10130.,0.0000,-5346.5,-7884.4,-487.04,-3436.9,-3581.5,-16063.,-1734.4,-1834.8,-5569.5,-3026.2,-6300.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
81.00000000000,0.12825E+06,9047.0,17382.,23129.,19863.,13410.,39366.,6764.6,18802.,3188.6,7869.9,9890.1,0.0000,-5339.6,-7879.5,-486.39,-3438.1,-3575.3,-16036.,-1734.4,-1827.4,-5567.5,-3027.1,-6295.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
82.00000000000,0.12622E+06,8990.4,17353.,22636.,19733.,12818.,38916.,6677.3,18617.,3158.7,7869.7,9712.2,0.0000,-5385.0,-7903.6,-490.15,-3439.7,-3603.9,-16009.,-1736.0,-1852.4,-5577.7,-3030.6,-6300.0,11092.,4957.8,3797.8,3564.4,6909.7,2381.0,8534.7,2466.3,3770.4,1125.4,1617.4,1948.3,0.0000,-14.708,-14.161,-1.7957,-12.272,-11.875,-50.235,-35.195,-3.5913,-31.939,-4.1438,-42.696
83.00000000000,0.12421E+06,8878.0,17334.,22002.,19366.,12555.,37834.,6617.2,18447.,3137.8,7794.7,9581.1,0.0000,-5352.9,-7901.7,-489.15,-3441.3,-3579.7,-15981.,-1735.6,-1830.1,-5568.0,-3029.9,-6290.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
84.00000000000,0.12026E+06,8797.6,17241.,21831.,18135.,12264.,37227.,6437.2,18287.,3051.7,7658.7,9445.1,0.0000,-5338.9,-7895.7,-487.79,-3442.7,-3571.2,-15955.,-1735.3,-1819.8,-5564.0,-3030.3,-6284.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
85.00000000000,0.11914E+06,8599.3,15082.,21488.,17055.,11992.,36547.,6303.2,17922.,2976.1,7540.8,9376.2,0.0000,-5326.8,-7888.4,-486.63,-3444.1,-3564.5,-15929.,-1735.1,-1812.0,-5561.5,-3030.9,-6279.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
86.00000000000,0.11546E+06,8389.3,14519.,21094.,16652.,11724.,36226.,6180.0,17642.,2948.4,7455.6,9266.9,0.0000,-5315.6,-7881.2,-485.59,-3445.5,-3558.5,-15903.,-1734.9,-1805.1,-5559.3,-3031.5,-6275.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
87.00000000000,0.11374E+06,8219.8,14441.,20747.,16318.,11427.,35455.,6098.8,17524.,2851.4,7276.7,9029.5,0.0000,-5305.1,-7874.4,-484.69,-3446.9,-3553.1,-15878.,-1734.8,-1798.6,-5557.3,-3032.1,-6270.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
88.00000000000,0.11265E+06,7977.2,14247.,20402.,15904.,11129.,34872.,5957.4,17208.,2793.4,7116.7,8875.5,0.0000,-5295.3,-7867.9,-483.87,-3448.3,-3548.1,-15854.,-1734.8,-1792.4,-5555.4,-3032.8,-6266.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
89.00000000000,0.11134E+06,7933.4,13929.,19956.,15765.,11082.,34200.,5735.1,16614.,2755.2,6863.4,8725.4,0.0000,-5286.0,-7861.5,-483.12,-3449.6,-3543.3,-15829.,-1734.8,-1786.5,-5553.6,-3033.4,-6262.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
90.00000000000,0.10907E+06,7732.0,13744.,19651.,15242.,11069.,33460.,5558.2,16206.,2741.0,6725.4,8637.2,0.0000,-5277.1,-7855.2,-482.42,-3451.0,-3538.7,-15805.,-1734.8,-1780.8,-5551.9,-3034.0,-6258.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
91.00000000000,0.10704E+06,7533.7,13632.,19369.,15030.,10908.,33102.,5271.5,16016.,2681.3,6612.3,8410.5,0.0000,-5268.6,-7849.3,-481.74,-3452.0,-3534.4,-15782.,-1734.8,-1775.4,-5550.1,-3034.6,-6254.6,70.849,31.668,24.259,22.768,44.136,15.209,54.516,15.754,24.084,7.1887,10.331,12.445,0.0000,-0.93052E-01,-0.90631E-01,-0.11470E-01,-0.78168E-01,-0.76186E-01,-0.31840,-0.22493,-0.22940E-01,-0.20395,-0.26622E-01,-0.27272
92.00000000000,0.10670E+06,7166.5,13508.,18991.,14866.,10770.,32561.,5115.9,15878.,2646.6,6508.8,8297.0,0.0000,-5260.3,-7843.7,-481.09,-3453.0,-3530.3,-15760.,-1734.8,-1770.3,-5548.3,-3035.2,-6250.4,173.10,77.374,59.271,55.628,107.84,37.160,133.20,38.491,58.843,17.564,25.243,30.406,0.0000,-0.22713,-0.22145,-0.28024E-01,-0.19093,-0.18624,-0.77723,-0.54958,-0.56048E-01,-0.49828,-0.65084E-01,-0.66633
93.00000000000,0.10656E+06,6880.5,13366.,18776.,14676.,10685.,32146.,5012.5,15661.,2611.6,6400.8,8151.5,0.0000,-5304.8,-7866.9,-484.82,-3454.3,-3555.7,-15740.,-1741.3,-1797.0,-5559.6,-3038.5,-6256.0,48135.,21516.,16482.,15468.,29986.,10333.,37039.,10703.,16363.,4884.1,7019.3,8455.1,0.0000,-63.243,-61.653,-7.7927,-53.155,-51.890,-215.93,-152.84,-15.585,-138.55,-18.112,-185.29
94.00000000000,0.10645E+06,6722.1,13323.,18659.,14611.,10409.,31734.,4962.1,15618.,2560.9,6274.8,8050.8,0.0000,-5272.3,-7863.5,-483.81,-3455.4,-3534.0,-15719.,-1739.8,-1776.8,-5550.6,-3037.5,-6247.5,760.86,340.09,260.52,244.51,473.98,163.33,585.46,169.18,258.64,77.201,110.95,133.65,0.0000,-0.99875,-0.97476,-0.12318,-0.83980,-0.82027,-3.4102,-2.4161,-0.24635,-2.1900,-0.28646,-2.9288
95.00000000000,0.10495E+06,6686.5,13282.,18446.,14493.,10307.,31494.,4789.6,15239.,2501.7,6128.2,7921.2,0.0000,-5259.3,-7855.6,-482.39,-3456.3,-3527.8,-15698.,-1738.4,-1768.2,-5546.9,-3037.5,-6242.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
96.00000000000,0.10460E+06,6584.6,13114.,18190.,14219.,10051.,31180.,4738.8,14820.,2475.4,6041.6,7793.3,0.0000,-5248.3,-7847.2,-481.14,-3457.2,-3523.2,-15679.,-1737.3,-1761.8,-5544.3,-3037.7,-6237.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
97.00000000000,0.10433E+06,6492.8,13050.,17919.,14031.,9791.3,30803.,4687.0,14635.,2459.1,5954.4,7662.4,0.0000,-5238.0,-7839.0,-480.08,-3458.1,-3519.1,-15660.,-1736.5,-1756.1,-5542.0,-3037.8,-6233.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
98.00000000000,0.10402E+06,6355.7,12933.,17595.,13931.,9611.9,30593.,4559.8,14613.,2367.2,5874.3,7539.7,0.0000,-5228.1,-7830.9,-479.15,-3458.9,-3515.0,-15641.,-1735.9,-1750.8,-5539.7,-3038.0,-6228.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
99.00000000000,0.10189E+06,6039.0,12712.,17474.,13533.,9398.6,30056.,4495.4,14441.,2333.7,5846.8,7446.2,0.0000,-5218.5,-7823.2,-478.32,-3459.7,-3510.7,-15623.,-1735.5,-1745.6,-5537.6,-3038.3,-6225.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
100.0000000000,99727.,5947.3,12609.,17189.,13250.,9229.7,29606.,4474.8,14126.,2321.4,5790.8,7384.0,0.0000,-5209.1,-7815.8,-477.56,-3460.4,-3506.5,-15605.,-1735.2,-1740.7,-5535.6,-3038.5,-6221.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
101.0000000000,98351.,5912.2,12520.,17124.,13094.,8993.4,29243.,4456.2,13925.,2284.4,5697.2,7298.8,0.0000,-5200.0,-7808.7,-476.84,-3461.2,-3502.4,-15588.,-1735.0,-1735.9,-5533.7,-3038.8,-6217.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
102.0000000000,97972.,5822.5,12524.,17099.,12896.,8866.9,29113.,4445.2,13830.,2213.1,5579.4,7191.0,0.0000,-5191.1,-7801.9,-476.16,-3461.9,-3498.3,-15571.,-1734.8,-1731.3,-5531.9,-3039.0,-6213.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
103.0000000000,96237.,5761.1,12528.,16690.,12736.,8899.3,28723.,4402.6,13790.,2129.1,5491.5,7119.0,0.0000,-5182.0,-7795.4,-475.50,-3462.6,-3494.4,-15552.,-1734.7,-1726.9,-5530.2,-3039.3,-6210.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
104.0000000000,95670.,5762.7,12498.,16340.,12441.,8849.5,28185.,4350.6,13482.,2093.7,5429.2,6945.4,0.0000,-5172.7,-7789.1,-474.84,-3463.3,-3490.4,-15529.,-1734.6,-1722.5,-5528.5,-3039.6,-6206.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
105.0000000000,94727.,5722.0,12480.,16219.,12303.,8830.4,27945.,4328.5,13258.,2069.6,5288.5,6737.1,0.0000,-5163.4,-7783.1,-474.17,-3463.9,-3486.6,-15508.,-1734.5,-1718.4,-5526.7,-3039.7,-6203.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
106.0000000000,89265.,5638.2,12453.,16053.,12214.,8687.0,27845.,4284.7,12792.,2023.8,5212.8,6627.3,0.0000,-5154.3,-7777.2,-473.49,-3464.5,-3482.9,-15487.,-1734.4,-1714.3,-5524.9,-3039.8,-6200.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
107.0000000000,84211.,5625.7,12440.,15941.,12073.,8566.6,27647.,4254.9,12463.,1980.4,5143.0,6532.3,0.0000,-5145.6,-7771.5,-472.81,-3465.1,-3479.2,-15467.,-1734.3,-1710.5,-5523.0,-3039.8,-6196.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
108.0000000000,81513.,5623.1,12446.,15783.,11996.,8508.8,27466.,4230.8,12250.,1962.7,5036.0,6446.8,0.0000,-5189.3,-7794.5,-476.49,-3466.1,-3504.1,-15449.,-1738.1,-1737.8,-5533.5,-3042.6,-6202.4,27755.,12406.,9503.4,8919.2,17290.,5958.1,21357.,6171.6,9434.9,2816.2,4047.4,4875.3,0.0000,-35.992,-35.559,-4.4933,-30.541,-29.969,-122.94,-88.187,-8.9866,-79.836,-10.522,-106.83
109.0000000000,81431.,5589.5,12418.,15386.,11927.,8334.4,27095.,4179.4,11849.,1952.2,4995.1,6365.3,0.0000,-5156.6,-7791.3,-475.44,-3466.8,-3483.1,-15431.,-1737.2,-1719.3,-5524.0,-3041.2,-6194.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
110.0000000000,80744.,5552.8,12392.,15114.,11867.,8259.1,26476.,4163.5,11739.,1912.7,4917.7,6214.3,0.0000,-5143.6,-7783.8,-473.98,-3467.4,-3477.4,-15413.,-1736.4,-1711.9,-5520.1,-3040.8,-6189.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
111.0000000000,79035.,5549.6,12259.,14987.,11816.,8115.4,26065.,4129.8,11592.,1863.8,4884.3,6099.8,0.0000,-5132.9,-7775.8,-472.68,-3467.9,-3473.2,-15396.,-1735.7,-1706.8,-5517.5,-3040.7,-6185.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
112.0000000000,77059.,5517.3,12237.,14605.,11657.,8078.8,25580.,4107.7,11432.,1835.9,4850.8,5968.8,0.0000,-5123.1,-7768.0,-471.57,-3468.4,-3469.4,-15380.,-1735.2,-1702.3,-5515.2,-3040.6,-6181.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
113.0000000000,74448.,5511.1,12239.,14178.,11436.,7968.2,24885.,4063.0,11397.,1825.5,4787.9,5869.1,0.0000,-5113.8,-7760.7,-470.60,-3468.9,-3465.7,-15364.,-1734.9,-1698.2,-5513.0,-3040.6,-6178.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
114.0000000000,73533.,5490.9,12191.,14131.,11127.,7961.9,24458.,4033.3,11254.,1814.3,4700.2,5744.3,0.0000,-5104.8,-7753.8,-469.73,-3469.3,-3462.2,-15349.,-1734.6,-1694.3,-5510.7,-3040.6,-6175.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
115.0000000000,72687.,5489.3,12104.,13914.,10990.,7866.9,24115.,3943.0,11216.,1804.4,4621.4,5693.5,0.0000,-5096.1,-7747.2,-468.94,-3469.7,-3458.7,-15335.,-1734.4,-1690.7,-5508.5,-3040.6,-6171.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
116.0000000000,71774.,5489.6,12083.,13675.,10804.,7814.8,23881.,3931.8,11112.,1802.6,4554.4,5609.2,0.0000,-5087.6,-7740.8,-468.19,-3470.1,-3455.4,-15320.,-1734.3,-1687.2,-5506.3,-3040.6,-6168.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
117.0000000000,70181.,5474.6,12064.,13528.,10389.,7639.1,23384.,3931.6,10717.,1793.4,4472.0,5597.6,0.0000,-5079.4,-7734.0,-467.47,-3470.4,-3452.0,-15306.,-1734.1,-1683.9,-5504.4,-3040.6,-6165.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
118.0000000000,70098.,5469.9,12055.,13514.,10077.,7635.4,23256.,3925.1,10493.,1781.0,4331.3,5556.0,0.0000,-5123.4,-7756.0,-471.03,-3471.0,-3477.3,-15293.,-1746.4,-1711.6,-5516.7,-3043.3,-6174.1,91278.,40800.,31254.,29333.,56862.,19594.,70236.,20296.,31028.,9261.6,13310.,16033.,0.0000,-117.39,-116.92,-14.777,-100.21,-98.342,-400.73,-290.12,-29.554,-262.42,-34.724,-351.30
119.0000000000,69055.,5345.5,11944.,13319.,9918.1,7622.8,23106.,3885.0,10303.,1765.6,4273.6,5502.9,0.0000,-5143.5,-7780.6,-474.25,-3471.8,-3485.1,-15280.,-1764.5,-1724.7,-5524.2,-3044.5,-6181.1,0.15574E+06,69615.,53327.,50049.,97022.,33433.,0.11984E+06,34631.,52942.,15803.,22711.,27357.,0.0000,-200.58,-199.74,-25.214,-171.14,-168.10,-683.16,-495.14,-50.427,-447.74,-59.272,-599.44
120.0000000000,68420.,5327.8,10376.,13061.,9798.8,7552.9,22757.,3863.7,10227.,1755.8,4224.9,5426.5,0.0000,-5107.1,-7775.2,-472.35,-3472.5,-3463.5,-15267.,-1756.7,-1702.5,-5514.5,-3042.6,-6174.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
121.0000000000,68105.,5305.3,10373.,12765.,9712.4,7507.0,22625.,3842.7,10175.,1751.4,4159.6,5378.7,0.0000,-5095.7,-7765.9,-470.25,-3473.6,-3458.9,-15256.,-1750.4,-1692.6,-5510.0,-3043.3,-6168.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
122.0000000000,67493.,5284.6,10375.,12541.,9651.3,7406.6,22479.,3799.9,10080.,1726.2,4109.8,5325.0,0.0000,-5137.3,-7785.9,-472.86,-3474.3,-3483.1,-15247.,-1753.7,-1716.3,-5520.5,-3046.7,-6173.4,58587.,26187.,20060.,18827.,36497.,12577.,45081.,13027.,19916.,5944.6,8543.4,10291.,0.0000,-75.484,-75.257,-9.4848,-64.418,-63.371,-256.53,-186.42,-18.970,-168.50,-22.348,-225.66
123.0000000000,67279.,5177.4,10313.,12375.,9601.2,7295.9,22124.,3802.4,10073.,1716.0,4030.2,5278.2,0.0000,-5103.9,-7778.5,-471.05,-3475.3,-3461.4,-15236.,-1748.3,-1695.2,-5510.2,-3045.3,-6164.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
124.0000000000,66947.,5125.0,10253.,12322.,9420.0,7255.5,21891.,3801.4,9865.6,1704.3,3992.4,5160.0,0.0000,-5089.3,-7766.9,-469.06,-3475.8,-3455.2,-15225.,-1744.2,-1685.8,-5505.7,-3045.7,-6157.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
125.0000000000,65271.,5125.5,10191.,12226.,9353.2,7147.2,21708.,3795.8,9670.2,1681.6,3979.0,5056.9,0.0000,-5077.9,-7754.5,-467.40,-3476.0,-3451.1,-15213.,-1741.3,-1679.0,-5502.0,-3045.6,-6153.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
126.0000000000,64523.,5114.6,10155.,12209.,9293.2,7134.4,21470.,3790.4,9644.2,1658.1,3909.9,5016.5,0.0000,-5067.7,-7743.2,-466.08,-3475.8,-3447.4,-15200.,-1739.1,-1673.2,-5498.8,-3045.9,-6148.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
127.0000000000,63189.,5048.1,10137.,12061.,9187.6,7121.2,21299.,3750.3,9520.0,1636.8,3864.6,4974.4,0.0000,-5057.7,-7734.9,-464.96,-3475.5,-3443.5,-15187.,-1737.7,-1668.2,-5496.4,-3046.6,-6144.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
128.0000000000,61716.,4995.9,10117.,12038.,9053.1,7093.6,20931.,3783.1,9414.2,1614.2,3835.8,4913.2,0.0000,-5048.3,-7725.9,-463.97,-3475.4,-3440.2,-15173.,-1736.6,-1663.7,-5494.6,-3047.3,-6140.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
129.0000000000,59924.,4963.3,10090.,11932.,8842.9,7095.6,20294.,3750.7,9307.4,1597.8,3777.1,4864.7,0.0000,-5039.3,-7716.1,-463.07,-3475.3,-3436.7,-15159.,-1735.8,-1659.4,-5492.6,-3048.1,-6137.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
130.0000000000,58043.,4970.1,10083.,11928.,8786.4,7101.0,19704.,3708.2,9261.6,1583.0,3731.1,4853.0,0.0000,-5082.7,-7735.2,-466.59,-3475.4,-3461.6,-15146.,-1739.4,-1686.0,-5503.1,-3051.0,-6143.1,29628.,13243.,10145.,9521.2,18457.,6360.2,22798.,6588.1,10072.,3006.2,4320.5,5204.3,0.0000,-37.905,-38.017,-4.7966,-32.506,-31.923,-128.88,-94.342,-9.5931,-85.209,-11.326,-114.16
131.0000000000,57047.,4930.4,10055.,11816.,8725.3,7078.4,19245.,3670.9,9081.0,1579.7,3673.3,4824.7,0.0000,-5101.9,-7757.1,-469.79,-3475.7,-3469.1,-15134.,-1743.0,-1698.7,-5506.4,-3052.5,-6144.4,36562.,16342.,12519.,11749.,22776.,7848.6,28133.,8129.7,12428.,3709.7,5331.5,6422.1,0.0000,-46.833,-46.962,-5.9190,-40.148,-39.452,-158.90,-116.43,-11.838,-105.14,-13.979,-140.88
132.0000000000,55652.,4930.1,10044.,11662.,8624.9,7004.7,18814.,3590.2,8995.2,1573.6,3623.2,4770.2,0.0000,-5064.3,-7748.6,-467.88,-3475.6,-3446.1,-15120.,-1740.7,-1676.3,-5495.2,-3050.9,-6135.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
133.0000000000,55365.,4909.1,10042.,11510.,8465.9,6841.1,18675.,3560.2,8923.6,1566.6,3574.3,4710.5,0.0000,-5048.7,-7735.6,-465.73,-3475.4,-3439.7,-15108.,-1738.8,-1666.7,-5490.7,-3050.6,-6129.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
134.0000000000,54763.,4866.5,10037.,11149.,8416.3,6705.7,18583.,3520.7,8845.5,1562.1,3523.2,4644.6,0.0000,-5036.7,-7722.9,-463.94,-3474.9,-3435.1,-15095.,-1737.3,-1659.6,-5487.6,-3050.3,-6125.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
135.0000000000,54108.,4830.8,9982.4,10831.,8420.1,6682.7,18536.,3504.8,8778.6,1551.7,3461.7,4520.5,0.0000,-5077.6,-7739.3,-466.83,-3474.6,-3459.6,-15085.,-1742.9,-1684.2,-5498.1,-3052.7,-6132.1,48263.,21573.,16525.,15510.,30066.,10361.,37137.,10732.,16406.,4897.1,7037.9,8477.5,0.0000,-61.666,-61.999,-7.8134,-52.945,-51.993,-209.10,-153.71,-15.627,-138.77,-18.463,-185.97
136.0000000000,54016.,4781.0,9908.1,10730.,8394.2,6662.0,18442.,3502.2,8685.3,1522.4,3444.6,4463.2,0.0000,-5042.8,-7730.9,-465.25,-3474.1,-3438.6,-15073.,-1740.5,-1664.0,-5488.6,-3050.8,-6124.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
137.0000000000,53759.,4788.0,9843.8,10662.,8395.1,6639.5,18232.,3501.3,8493.6,1496.7,3398.8,4456.9,0.0000,-5028.5,-7719.0,-463.42,-3473.5,-3432.6,-15062.,-1738.6,-1655.0,-5484.7,-3050.3,-6119.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
138.0000000000,53190.,4787.6,9216.1,10606.,8395.7,6638.2,18056.,3472.9,8442.3,1473.5,3339.6,4421.4,0.0000,-5016.8,-7707.6,-461.84,-3472.7,-3428.0,-15052.,-1737.2,-1648.3,-5482.1,-3050.1,-6115.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
139.0000000000,52747.,4773.7,8248.9,10499.,8392.4,6621.2,17902.,3426.6,8360.6,1445.7,3317.6,4366.6,0.0000,-5006.0,-7696.7,-460.52,-3472.0,-3424.0,-15042.,-1736.1,-1642.6,-5480.2,-3049.9,-6111.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
140.0000000000,52198.,4775.6,8252.9,10382.,8296.4,6521.0,17600.,3389.6,8338.4,1438.5,3281.7,4290.1,0.0000,-4996.2,-7686.5,-459.38,-3471.3,-3420.1,-15032.,-1735.3,-1637.4,-5478.6,-3049.8,-6108.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
141.0000000000,52060.,4775.2,8230.3,10090.,8203.1,6517.9,17330.,3334.1,8306.3,1437.8,3241.6,4240.4,0.0000,-4986.9,-7677.1,-458.37,-3470.6,-3416.3,-15022.,-1734.8,-1632.6,-5477.0,-3049.4,-6105.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
142.0000000000,50583.,4733.0,8197.2,9901.7,8207.5,6415.1,17078.,3318.2,8204.6,1422.2,3209.0,4204.5,0.0000,-4977.8,-7668.6,-457.46,-3469.9,-3412.5,-15013.,-1734.4,-1628.1,-5475.6,-3049.2,-6102.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
143.0000000000,50053.,4710.6,8147.7,9838.6,8226.3,6307.1,16858.,3282.5,8083.8,1403.2,3175.8,4197.6,0.0000,-4969.0,-7660.6,-456.61,-3469.4,-3408.6,-15004.,-1734.1,-1623.9,-5474.2,-3048.8,-6099.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
144.0000000000,49737.,4714.4,8133.5,9787.0,8190.9,6253.2,16736.,3254.5,8083.2,1399.8,3166.9,4196.6,0.0000,-5012.2,-7680.5,-460.14,-3469.1,-3433.1,-14995.,-1748.6,-1650.3,-5487.7,-3051.1,-6108.5,0.10892E+06,48684.,37293.,35001.,67851.,23381.,83809.,24219.,37024.,11051.,15883.,19132.,0.0000,-138.13,-139.68,-17.633,-119.05,-116.72,-468.73,-347.04,-35.266,-313.13,-41.721,-419.73
145.0000000000,49218.,4715.5,8131.5,9702.6,8194.3,6141.9,16507.,3213.0,8078.0,1389.4,3099.9,4180.9,0.0000,-5031.3,-7702.4,-463.33,-3468.9,-3440.4,-14987.,-1746.1,-1663.0,-5491.7,-3051.7,-6110.9,8943.5,3997.6,3062.3,2874.0,5571.4,1919.9,6881.7,1988.7,3040.2,907.45,1304.2,1570.9,0.0000,-11.357,-11.482,-1.4479,-9.7830,-9.5982,-38.455,-28.498,-2.8957,-25.712,-3.4265,-34.465
146.0000000000,48674.,4717.7,8066.8,9508.3,8200.2,6054.9,16358.,3167.7,8034.4,1385.7,3089.6,4141.4,0.0000,-5046.0,-7722.5,-465.73,-3468.9,-3445.6,-14978.,-1765.8,-1671.9,-5496.9,-3052.2,-6116.1,0.16999E+06,75982.,58204.,54627.,0.10590E+06,36491.,0.13080E+06,37799.,57785.,17248.,24788.,29859.,0.0000,-216.15,-218.48,-27.520,-186.06,-182.66,-730.30,-541.79,-55.040,-488.73,-65.139,-655.12
147.0000000000,48418.,4736.1,8055.0,9343.0,8215.1,6018.9,16323.,3142.3,7978.7,1376.2,3080.7,4150.2,0.0000,-5008.5,-7712.5,-463.21,-3469.2,-3423.9,-14969.,-1757.4,-1648.3,-5486.8,-3050.5,-6108.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
148.0000000000,47999.,4750.5,8086.8,9281.8,8202.8,5993.4,16298.,3117.8,7950.6,1363.7,3068.8,4136.4,0.0000,-4995.9,-7702.8,-460.64,-3469.4,-3418.2,-14965.,-1750.8,-1638.4,-5483.2,-3052.1,-6103.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
149.0000000000,47664.,4715.1,8067.6,9269.9,8157.1,5966.5,15994.,3077.5,7825.0,1353.8,3049.9,4103.6,0.0000,-5036.8,-7717.6,-462.87,-3470.4,-3441.8,-14958.,-1749.1,-1662.2,-5492.8,-3056.3,-6107.4,23746.,10614.,8130.6,7630.9,14793.,5097.5,18272.,5280.1,8072.0,2409.4,3462.7,4171.0,0.0000,-30.217,-30.557,-3.8443,-25.992,-25.549,-101.88,-75.752,-7.6885,-68.339,-9.1223,-91.590
150.0000000000,47042.,4702.6,8066.7,9260.6,8104.3,5874.2,15843.,3052.8,7679.9,1351.1,3029.7,4042.9,0.0000,-5001.8,-7707.4,-460.88,-3469.9,-3419.5,-14951.,-1744.7,-1641.9,-5481.9,-3056.7,-6098.2,185.18,82.772,63.406,59.509,115.36,39.752,142.49,41.176,62.949,18.789,27.004,32.527,0.0000,-0.23534,-0.23822,-0.29979E-01,-0.20251,-0.19890,-0.79378,-0.59080,-0.59958E-01,-0.53299,-0.71155E-01,-0.71428
151.0000000000,46650.,4664.9,8017.2,9154.4,7988.5,5836.8,15633.,3027.4,7625.5,1347.1,3024.1,3958.6,0.0000,-4986.1,-7695.1,-458.76,-3469.1,-3413.3,-14943.,-1741.5,-1633.2,-5477.4,-3058.8,-6092.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
152.0000000000,46461.,4617.9,8020.2,8985.3,7946.9,5727.6,15564.,3009.3,7619.2,1343.1,3003.1,3944.1,0.0000,-4974.1,-7683.1,-456.99,-3468.0,-3408.5,-14936.,-1739.2,-1627.0,-5473.9,-3061.1,-6088.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
153.0000000000,46257.,4579.9,8018.8,8768.0,7936.3,5450.9,15530.,3003.6,7608.9,1340.5,2987.9,3917.2,0.0000,-4963.3,-7671.8,-455.54,-3466.6,-3404.3,-14929.,-1737.5,-1621.8,-5471.2,-3062.1,-6085.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
154.0000000000,45071.,4578.3,8005.0,8480.3,7898.9,5433.7,15279.,2958.1,7599.7,1329.0,2985.3,3873.2,0.0000,-5005.3,-7689.5,-458.61,-3465.7,-3428.8,-14923.,-1736.9,-1647.6,-5480.6,-3065.4,-6090.1,3557.4,1590.1,1218.1,1143.2,2216.1,763.67,2737.3,791.02,1209.3,360.96,518.76,624.87,0.0000,-4.5075,-4.5737,-0.57592,-3.8849,-3.8119,-15.200,-11.351,-1.1518,-10.240,-1.3673,-13.723
155.0000000000,44259.,4532.5,7969.2,8429.0,7875.2,5375.1,15153.,2878.7,7599.0,1299.7,2942.1,3852.9,0.0000,-4972.1,-7681.2,-457.13,-3464.5,-3407.5,-14916.,-1736.0,-1629.2,-5470.5,-3063.5,-6081.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
156.0000000000,44043.,4504.9,7478.3,8346.0,7856.0,5141.0,14901.,2853.7,7497.2,1286.6,2896.4,3811.1,0.0000,-4959.0,-7669.3,-455.32,-3463.1,-3401.2,-14910.,-1735.3,-1621.5,-5466.8,-3062.2,-6077.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
157.0000000000,43742.,4476.9,6275.3,8272.7,7890.4,5067.7,14653.,2796.4,7354.9,1264.6,2858.0,3801.1,0.0000,-4948.7,-7657.5,-453.75,-3461.7,-3396.5,-14903.,-1734.8,-1616.1,-5464.8,-3060.5,-6074.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
158.0000000000,43034.,4398.2,6259.1,8251.7,7899.9,5056.0,14616.,2761.2,7334.3,1256.5,2839.3,3777.6,0.0000,-4938.2,-7647.4,-452.41,-3459.8,-3392.4,-14897.,-1734.5,-1611.6,-5463.3,-3059.1,-6072.4,913.02,408.10,312.62,293.40,568.77,196.00,702.54,203.02,310.36,92.640,133.14,160.37,0.0000,-1.1514,-1.1724,-0.14781,-0.99407,-0.97351,-3.8896,-2.9132,-0.29562,-2.6280,-0.35082,-3.5219
159.0000000000,42752.,4383.3,6223.8,8251.1,7254.6,5055.3,14526.,2720.8,7264.5,1238.4,2839.2,3743.6,0.0000,-4979.8,-7665.9,-455.55,-3458.1,-3417.3,-14891.,-1739.4,-1637.8,-5474.9,-3060.6,-6079.8,38409.,17168.,13151.,12343.,23927.,8245.2,29555.,8540.5,13056.,3897.2,5600.9,6746.6,0.0000,-48.494,-49.356,-6.2181,-41.855,-41.026,-163.50,-122.55,-12.436,-110.55,-14.760,-148.19
160.0000000000,42355.,4330.5,6158.6,8140.3,7234.0,4903.5,14351.,2677.5,7196.7,1220.1,2832.4,3701.6,0.0000,-4946.1,-7658.8,-454.13,-3456.4,-3396.5,-14883.,-1737.9,-1619.9,-5466.4,-3058.9,-6073.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
161.0000000000,42173.,4328.6,6163.1,8128.8,7195.1,4885.5,14068.,2673.7,7095.1,1179.7,2817.5,3639.9,0.0000,-4931.7,-7648.1,-452.38,-3454.5,-3390.9,-14876.,-1736.7,-1612.5,-5463.2,-3059.2,-6069.5,129.61,57.935,44.380,41.652,80.744,27.824,99.734,28.821,44.060,13.151,18.901,22.767,0.0000,-0.16329,-0.16649,-0.20983E-01,-0.14104,-0.13814,-0.55099,-0.41356,-0.41967E-01,-0.37304,-0.49815E-01,-0.50025
162.0000000000,41944.,4317.3,6132.6,8040.8,7147.4,4759.2,13896.,2669.3,6998.5,1144.2,2801.4,3583.8,0.0000,-4920.2,-7638.1,-450.85,-3452.5,-3386.6,-14869.,-1735.7,-1607.5,-5461.5,-3059.8,-6066.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
163.0000000000,41711.,4319.9,6130.8,8037.2,7159.4,4696.3,13889.,2588.5,6906.3,1142.1,2779.8,3546.4,0.0000,-4910.2,-7628.8,-449.55,-3450.3,-3382.8,-14862.,-1734.9,-1603.8,-5460.1,-3060.0,-6064.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
164.0000000000,41415.,4308.6,6104.7,7922.2,7195.8,4667.7,13601.,2493.1,6820.0,1132.9,2758.6,3509.7,0.0000,-4901.3,-7620.0,-448.41,-3448.8,-3379.4,-14856.,-1734.4,-1600.4,-5458.9,-3059.3,-6061.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
165.0000000000,41326.,4309.2,6082.3,7903.8,7210.1,4629.1,13542.,2439.6,6660.1,1131.6,2714.6,3464.0,0.0000,-4944.4,-7639.0,-451.71,-3447.7,-3404.6,-14851.,-1737.4,-1627.1,-5470.3,-3061.3,-6068.0,24421.,10916.,8361.7,7847.7,15213.,5242.4,18791.,5430.2,8301.4,2477.9,3561.1,4289.6,0.0000,-30.705,-31.357,-3.9535,-26.550,-25.993,-103.56,-77.916,-7.9071,-70.280,-9.3891,-94.326
166.0000000000,41123.,4296.2,6044.7,7868.5,7157.4,4627.5,13485.,2388.3,6598.4,1129.0,2705.6,3424.3,0.0000,-4963.5,-7661.7,-454.74,-3446.7,-3412.0,-14846.,-1765.9,-1639.8,-5479.5,-3062.1,-6076.7,0.21818E+06,97522.,74705.,70113.,0.13592E+06,46836.,0.16788E+06,48514.,74166.,22138.,31816.,38324.,0.0000,-274.72,-280.43,-35.321,-237.38,-232.54,-924.61,-696.29,-70.643,-627.89,-83.895,-842.92
167.0000000000,41013.,4273.8,6045.1,7817.3,7032.7,4654.8,13341.,2336.6,6480.9,1128.1,2689.6,3407.7,0.0000,-4979.0,-7684.3,-457.07,-3446.0,-3419.9,-14840.,-1760.0,-1649.0,-5482.9,-3062.7,-6080.0,16276.,7275.1,5572.9,5230.4,10139.,3493.9,12524.,3619.1,5532.7,1651.5,2373.4,2858.9,0.0000,-20.531,-20.948,-2.6350,-17.727,-17.391,-68.962,-51.955,-5.2699,-46.847,-6.2597,-62.916
168.0000000000,40943.,4262.8,6023.7,7799.4,7004.2,4624.8,13268.,2269.4,6380.5,1129.7,2694.4,3378.6,0.0000,-4943.9,-7679.1,-454.52,-3445.7,-3397.9,-14838.,-1752.8,-1625.9,-5471.4,-3062.7,-6070.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
169.0000000000,40857.,4260.8,5974.2,7737.7,7007.3,4615.2,13024.,2178.7,6393.7,1118.5,2663.7,3340.4,0.0000,-4980.2,-7694.3,-456.24,-3445.8,-3419.8,-14835.,-1749.5,-1646.8,-5479.5,-3065.5,-6073.7,16210.,7245.4,5550.2,5209.0,10098.,3479.7,12473.,3604.3,5510.1,1644.7,2363.7,2847.2,0.0000,-20.474,-20.887,-2.6242,-17.658,-17.329,-68.642,-51.768,-5.2484,-46.686,-6.2452,-62.748
170.0000000000,40775.,4201.3,5917.3,7567.4,7012.1,4494.0,12982.,2128.5,6360.2,1115.1,2663.8,3313.6,0.0000,-4995.1,-7709.4,-458.10,-3444.7,-3425.2,-14831.,-1745.6,-1656.5,-5480.0,-3068.2,-6072.4,4773.0,2133.4,1634.3,1533.8,2973.3,1024.6,3672.6,1061.3,1622.5,484.29,696.01,838.38,0.0000,-6.0339,-6.1549,-0.77270,-5.2020,-5.1068,-20.198,-15.244,-1.5454,-13.749,-1.8393,-18.483
171.0000000000,40776.,4141.6,5890.5,7421.2,6989.7,4379.3,12831.,2119.3,6321.3,1088.6,2623.4,3295.0,0.0000,-4954.3,-7694.5,-455.31,-3442.8,-3400.7,-14825.,-1742.1,-1632.6,-5467.0,-3066.1,-6061.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
172.0000000000,40754.,4024.2,5862.1,7231.2,6959.5,4365.9,12618.,2085.0,6298.2,1069.4,2616.1,3264.5,0.0000,-4936.0,-7677.2,-452.59,-3440.6,-3393.3,-14819.,-1739.6,-1622.3,-5461.3,-3065.8,-6056.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
173.0000000000,40558.,3975.0,5855.4,7205.5,6937.6,4364.8,12524.,2040.3,6260.8,1068.0,2594.7,3223.8,0.0000,-4921.3,-7662.1,-450.42,-3438.3,-3388.1,-14815.,-1737.8,-1615.4,-5458.1,-3065.8,-6052.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
174.0000000000,40505.,3940.2,5823.6,7207.6,6937.7,4245.9,12379.,2012.2,6223.0,1052.0,2572.6,3214.7,0.0000,-4908.2,-7647.7,-448.68,-3436.0,-3383.5,-14810.,-1736.5,-1609.7,-5455.8,-3066.2,-6048.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
175.0000000000,40462.,3919.5,5786.0,7209.0,6903.9,4174.4,12315.,1972.3,6212.8,1037.4,2531.4,3158.7,0.0000,-4896.2,-7634.3,-447.25,-3433.9,-3379.1,-14805.,-1735.6,-1604.7,-5453.7,-3066.4,-6045.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
176.0000000000,40276.,3908.6,5723.4,7210.6,6897.9,4165.3,12255.,1918.6,6168.2,1015.2,2509.8,3132.4,0.0000,-4885.4,-7622.2,-446.03,-3431.9,-3374.9,-14800.,-1735.0,-1600.1,-5451.9,-3066.0,-6042.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
177.0000000000,39763.,3905.1,5723.2,7173.1,6892.9,4135.3,12209.,1867.6,5963.9,1009.9,2497.2,3081.8,0.0000,-4874.9,-7610.7,-444.96,-3430.0,-3371.0,-14796.,-1734.5,-1595.9,-5450.2,-3065.2,-6040.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
178.0000000000,39696.,3905.7,5708.3,7073.0,6802.1,3963.9,12131.,1850.0,5849.0,999.34,2490.2,3065.4,0.0000,-4864.7,-7600.4,-444.00,-3428.2,-3367.1,-14791.,-1734.1,-1592.1,-5448.7,-3064.6,-6037.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
179.0000000000,39625.,3840.5,5705.5,7043.6,6795.9,3874.1,11984.,1851.6,5845.4,997.04,2481.6,3038.3,0.0000,-4854.9,-7591.1,-443.10,-3426.4,-3363.3,-14787.,-1733.9,-1588.7,-5447.8,-3064.2,-6035.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
180.0000000000,39565.,3761.5,5683.7,6993.3,6831.4,3864.0,11884.,1827.7,5844.2,995.24,2454.3,3006.0,0.0000,-4845.5,-7583.0,-442.26,-3424.8,-3359.6,-14782.,-1733.7,-1585.5,-5446.4,-3063.8,-6033.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
181.0000000000,39559.,3715.3,5668.4,6940.4,6777.4,3880.0,11779.,1806.3,5820.0,968.40,2437.0,2989.1,0.0000,-4887.5,-7602.3,-445.76,-3423.6,-3384.6,-14779.,-1740.9,-1612.3,-5458.4,-3066.1,-6041.5,54108.,24185.,18526.,17388.,33707.,11615.,41634.,12031.,18393.,5490.1,7890.2,9504.1,0.0000,-67.567,-69.484,-8.7596,-58.603,-57.205,-227.45,-172.80,-17.519,-155.83,-20.852,-209.98
182.0000000000,39533.,3706.9,5656.9,6925.4,6769.7,3830.4,11748.,1742.7,5796.3,947.93,2415.2,2966.7,0.0000,-4854.6,-7596.7,-444.63,-3422.4,-3363.6,-14774.,-1739.1,-1595.7,-5450.1,-3064.9,-6035.1,574.70,256.88,196.78,184.68,358.01,123.37,442.21,127.79,195.36,58.312,83.804,100.95,0.0000,-0.71689,-0.73789,-0.93038E-01,-0.62199,-0.60674,-2.4144,-1.8353,-0.18608,-1.6551,-0.22147,-2.2306
183.0000000000,39490.,3708.3,5640.2,6903.5,6784.5,3759.5,11761.,1722.7,5808.4,940.54,2391.8,2962.3,0.0000,-4892.6,-7615.8,-447.39,-3421.3,-3386.4,-14770.,-1739.1,-1619.3,-5459.1,-3067.0,-6040.4,12127.,5420.6,4152.3,3897.1,7554.7,2603.3,9331.4,2696.6,4122.4,1230.5,1768.4,2130.2,0.0000,-15.146,-15.583,-1.9633,-13.136,-12.821,-50.919,-38.727,-3.9265,-34.924,-4.6742,-47.077
184.0000000000,39419.,3699.7,5624.9,6865.6,6771.8,3706.5,11751.,1697.4,5799.0,936.15,2362.9,2949.9,0.0000,-4858.0,-7609.2,-445.68,-3420.2,-3364.9,-14765.,-1737.5,-1601.3,-5449.4,-3064.8,-6032.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
185.0000000000,39380.,3630.3,5620.1,6802.3,6763.9,3682.8,11693.,1696.7,5709.0,934.54,2357.6,2930.7,0.0000,-4843.9,-7598.7,-443.73,-3419.2,-3358.9,-14761.,-1736.2,-1593.9,-5445.7,-3063.9,-6028.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
186.0000000000,39335.,3588.9,5602.8,6686.8,6696.6,3638.4,11624.,1694.1,5677.7,935.62,2356.0,2924.1,0.0000,-4832.1,-7587.9,-442.08,-3418.0,-3354.4,-14756.,-1735.3,-1588.9,-5444.1,-3063.4,-6025.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
187.0000000000,39261.,3552.9,5579.8,6671.2,6673.1,3621.6,11506.,1685.8,5677.0,932.00,2347.4,2922.8,0.0000,-4821.5,-7577.6,-440.72,-3416.6,-3350.5,-14752.,-1734.6,-1584.8,-5442.3,-3062.9,-6022.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
188.0000000000,39259.,3492.7,5554.6,6671.6,6648.3,3590.7,11443.,1679.0,5662.4,917.84,2345.8,2924.1,0.0000,-4811.5,-7568.8,-439.56,-3415.5,-3347.0,-14747.,-1734.1,-1581.1,-5440.9,-3062.5,-6020.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
189.0000000000,39253.,3438.2,5485.8,6667.8,6635.7,3557.8,11386.,1677.5,5629.5,892.61,2343.1,2918.5,0.0000,-4802.0,-7559.6,-438.55,-3414.4,-3343.7,-14742.,-1733.7,-1577.8,-5439.8,-3062.3,-6018.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
190.0000000000,39257.,3396.0,5387.1,6660.9,6621.4,3538.6,11328.,1665.6,5611.3,859.16,2307.5,2915.1,0.0000,-4793.0,-7550.9,-437.65,-3413.2,-3340.1,-14738.,-1733.4,-1574.8,-5438.9,-3062.4,-6016.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
191.0000000000,39225.,3333.1,5353.2,6629.6,6556.9,3485.1,11317.,1621.7,5614.2,833.49,2287.2,2905.8,0.0000,-4784.4,-7543.1,-436.81,-3411.9,-3336.6,-14734.,-1733.2,-1572.0,-5438.0,-3062.4,-6014.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
192.0000000000,39220.,3292.8,5309.6,6573.2,6563.0,3479.0,11206.,1609.7,5596.8,828.46,2272.2,2892.3,0.0000,-4775.8,-7535.9,-436.02,-3410.6,-3333.2,-14730.,-1733.1,-1569.5,-5437.2,-3062.3,-6012.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
193.0000000000,38617.,3280.5,5294.4,6570.8,6566.0,3476.3,11078.,1602.3,5515.5,824.13,2265.1,2845.7,0.0000,-4767.3,-7528.7,-435.27,-3409.3,-3330.0,-14755.,-1732.9,-1567.1,-5436.5,-3062.0,-6010.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
194.0000000000,38603.,3237.1,5296.0,6543.3,6568.9,3476.9,10965.,1596.9,5516.7,815.72,2252.6,2830.3,0.0000,-4759.1,-7521.7,-434.55,-3408.2,-3326.7,-14751.,-1732.8,-1564.8,-5435.6,-3061.7,-6008.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
195.0000000000,38568.,3165.7,5294.9,6531.5,6568.4,3479.7,10899.,1596.1,5483.8,812.17,2252.7,2830.7,0.0000,-4751.2,-7515.1,-433.85,-3407.0,-3323.4,-14745.,-1732.7,-1562.6,-5434.7,-3061.4,-6006.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
196.0000000000,38557.,3104.5,5299.4,6538.5,6528.5,3496.0,10856.,1565.6,5388.4,810.22,2252.8,2824.0,0.0000,-4794.6,-7536.2,-437.45,-3406.2,-3348.6,-14739.,-1734.5,-1589.8,-5445.8,-3064.1,-6013.1,13707.,6126.6,4693.2,4404.7,8538.7,2942.4,10547.,3047.8,4659.3,1390.8,1998.8,2407.6,0.0000,-16.919,-17.534,-2.2190,-14.757,-14.312,-57.148,-43.753,-4.4380,-39.458,-5.2865,-53.311
197.0000000000,38560.,3079.5,5259.2,6540.9,6463.5,3449.0,10778.,1563.8,5393.3,808.11,2245.2,2805.8,0.0000,-4814.2,-7560.1,-440.74,-3405.4,-3356.4,-14733.,-1753.4,-1603.9,-5452.9,-3065.3,-6019.5,0.14224E+06,63580.,48704.,45711.,88612.,30535.,0.10945E+06,31629.,48353.,14433.,20742.,24985.,0.0000,-175.84,-182.14,-23.028,-153.27,-148.71,-592.75,-454.11,-46.056,-409.47,-54.872,-553.34
198.0000000000,38559.,3072.2,5188.4,6545.6,6449.1,3402.7,10663.,1561.1,5302.5,801.64,2236.3,2797.5,0.0000,-4829.5,-7582.3,-443.26,-3404.6,-3361.9,-14728.,-1758.5,-1614.1,-5457.7,-3066.0,-6024.3,75081.,33560.,25708.,24127.,46772.,16117.,57772.,16695.,25522.,7618.1,10949.,13188.,0.0000,-92.943,-96.237,-12.155,-80.951,-78.573,-312.72,-239.71,-24.310,-216.13,-28.967,-292.12
199.0000000000,38561.,3083.5,5146.4,6550.9,6456.6,3397.0,10642.,1560.0,5259.9,789.22,2222.8,2777.6,0.0000,-4842.9,-7602.0,-445.17,-3404.0,-3367.4,-14723.,-1753.6,-1622.6,-5459.0,-3066.4,-6025.3,14003.,6259.2,4794.7,4500.0,8723.4,3006.0,10775.,3113.7,4760.1,1420.8,2042.0,2459.7,0.0000,-17.360,-17.969,-2.2670,-15.109,-14.677,-58.304,-44.713,-4.5340,-40.311,-5.4034,-54.501
200.0000000000,38515.,3079.2,5122.9,6532.1,6430.8,3373.6,10681.,1563.9,5202.4,795.99,2230.1,2775.0,0.0000,-4857.4,-7620.2,-446.69,-3404.0,-3373.2,-14719.,-1751.0,-1629.9,-5459.1,-3067.6,-6024.3,22722.,10157.,7780.2,7301.9,14155.,4877.8,17484.,5052.5,7724.1,2305.5,3313.5,3991.2,0.0000,-28.234,-29.200,-3.6786,-24.542,-23.857,-94.613,-72.572,-7.3571,-65.433,-8.7771,-88.491
201.0000000000,38273.,3022.0,5083.4,6510.1,6389.6,3346.0,10666.,1545.5,5146.0,789.14,2215.9,2763.6,0.0000,-4818.1,-7610.3,-443.60,-3403.1,-3348.9,-14716.,-1745.9,-1605.9,-5447.2,-3066.2,-6013.7,345.48,154.42,118.29,111.02,215.22,74.163,265.83,76.820,117.44,35.054,50.379,60.684,0.0000,-0.42884,-0.44387,-0.55930E-01,-0.37276,-0.36206,-1.4381,-1.1035,-0.11186,-0.99502,-0.13350,-1.3460
202.0000000000,38246.,3023.9,5070.0,6491.2,6331.1,3353.6,10629.,1536.5,5127.6,787.31,2199.3,2770.5,0.0000,-4852.5,-7621.8,-444.94,-3403.0,-3369.7,-14712.,-1742.7,-1625.8,-5454.4,-3068.7,-6016.2,3784.4,1691.6,1295.8,1216.1,2357.5,812.39,2912.0,841.49,1286.4,383.99,551.86,664.74,0.0000,-4.7020,-4.8649,-0.61266,-4.0856,-3.9697,-15.745,-12.089,-1.2253,-10.900,-1.4626,-14.749
203.0000000000,38060.,2991.9,5063.9,6480.7,6290.1,3354.4,10607.,1533.7,5135.3,787.43,2183.3,2768.3,0.0000,-4866.4,-7635.2,-446.55,-3402.3,-3375.3,-14708.,-1740.7,-1634.9,-5455.3,-3070.1,-6015.3,6003.7,2683.5,2055.7,1929.3,3740.0,1288.8,4619.7,1335.0,2040.8,609.17,875.48,1054.6,0.0000,-7.4666,-7.7232,-0.97195,-6.4843,-6.3021,-24.965,-19.179,-1.9439,-17.293,-2.3208,-23.403
204.0000000000,37618.,2900.2,5063.5,6472.1,6293.1,3337.1,10551.,1538.1,5121.9,782.14,2177.0,2761.4,0.0000,-4825.6,-7620.2,-443.64,-3401.1,-3351.1,-14702.,-1738.4,-1610.7,-5442.9,-3068.1,-6005.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
205.0000000000,37584.,2839.4,5029.7,6433.2,6292.1,3333.2,10463.,1539.9,5074.3,779.21,2186.2,2755.2,0.0000,-4807.5,-7603.4,-440.83,-3399.6,-3343.5,-14698.,-1736.8,-1600.0,-5438.4,-3068.2,-6000.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
206.0000000000,37586.,2826.8,5022.7,6427.8,6311.1,3313.1,10413.,1535.2,5085.6,773.62,2186.8,2740.6,0.0000,-4792.9,-7587.1,-438.60,-3397.8,-3338.1,-14693.,-1735.6,-1592.7,-5436.1,-3068.6,-5997.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
207.0000000000,37432.,2790.5,5017.9,6428.7,6288.6,3337.1,10420.,1524.6,5067.8,769.42,2190.6,2724.2,0.0000,-4780.0,-7572.0,-436.84,-3396.1,-3333.1,-14689.,-1734.7,-1586.6,-5434.3,-3069.1,-5994.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
208.0000000000,37390.,2781.8,5024.1,6421.7,6254.2,3330.2,10426.,1514.9,5059.8,763.43,2189.0,2710.0,0.0000,-4819.7,-7586.0,-439.53,-3394.7,-3357.0,-14687.,-1735.0,-1611.3,-5444.4,-3072.3,-6000.6,6306.8,2819.0,2159.4,2026.7,3928.8,1353.9,4852.9,1402.4,2143.9,639.92,919.67,1107.8,0.0000,-7.8066,-8.0978,-1.0210,-6.7929,-6.5821,-26.160,-20.157,-2.0420,-18.167,-2.4386,-24.606
209.0000000000,36905.,2754.1,5019.1,6363.1,6254.4,3288.3,10432.,1511.3,5051.9,761.60,2182.9,2699.5,0.0000,-4785.1,-7575.5,-437.73,-3393.2,-3335.2,-14683.,-1734.3,-1592.6,-5435.1,-3070.7,-5993.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
210.0000000000,36552.,2752.5,4959.2,6332.8,6250.6,3297.7,10448.,1508.3,5045.9,758.69,2171.0,2686.5,0.0000,-4821.6,-7589.5,-439.96,-3391.9,-3357.0,-14680.,-1736.7,-1614.6,-5443.9,-3072.8,-5998.8,21072.,9418.7,7215.0,6771.5,13127.,4523.4,16214.,4685.5,7163.0,2138.1,3072.8,3701.3,0.0000,-26.078,-27.061,-3.4113,-22.692,-21.974,-87.318,-67.358,-6.8227,-60.694,-8.1482,-82.231
211.0000000000,36470.,2747.3,4897.6,6248.6,6253.8,3286.9,10430.,1502.3,4999.4,757.00,2158.4,2665.5,0.0000,-4785.5,-7578.3,-437.82,-3390.4,-3334.7,-14676.,-1735.6,-1594.9,-5434.3,-3070.7,-5991.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
212.0000000000,36423.,2759.7,4847.5,6168.5,6217.1,3278.5,10435.,1496.1,4987.7,754.78,2155.3,2650.6,0.0000,-4769.7,-7563.4,-435.52,-3388.7,-3327.8,-14672.,-1734.7,-1586.6,-5431.0,-3069.7,-5987.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
213.0000000000,36384.,2754.2,4809.3,6148.5,6175.5,3221.0,10335.,1486.9,4900.7,752.19,2153.1,2634.4,0.0000,-4757.0,-7549.1,-433.58,-3386.9,-3322.7,-14669.,-1734.0,-1580.8,-5429.3,-3069.2,-5985.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
214.0000000000,36343.,2720.8,4807.4,6150.2,5593.6,3209.0,10330.,1481.8,4844.5,751.13,2149.4,2616.2,0.0000,-4745.8,-7536.2,-431.95,-3385.2,-3318.0,-14665.,-1733.5,-1576.0,-5428.0,-3068.6,-5983.0,313.47,140.12,107.33,100.74,195.28,67.292,241.21,69.703,106.56,31.806,45.711,55.062,0.0000,-0.38591,-0.40166,-0.50748E-01,-0.33650,-0.32480,-1.2965,-1.0022,-0.10150,-0.90274,-0.12118,-1.2238
215.0000000000,36304.,2703.4,4760.1,6134.1,5571.7,3187.5,10295.,1479.3,4820.5,747.77,2147.4,2595.7,0.0000,-4735.2,-7524.5,-430.55,-3383.6,-3313.7,-14662.,-1733.1,-1571.8,-5426.9,-3068.0,-5981.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
216.0000000000,36300.,2630.6,4692.4,6119.3,5569.6,3174.3,10261.,1476.8,4809.1,745.86,2143.6,2580.8,0.0000,-4724.9,-7513.7,-429.31,-3382.0,-3309.6,-14658.,-1732.7,-1568.0,-5425.7,-3067.4,-5979.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
217.0000000000,36301.,2552.3,4647.5,6097.9,5548.0,3153.0,10250.,1470.6,4805.2,744.64,2134.7,2586.6,0.0000,-4715.0,-7503.5,-428.19,-3380.4,-3305.6,-14654.,-1732.5,-1564.5,-5424.7,-3066.7,-5977.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
218.0000000000,36310.,2545.5,4475.4,6086.5,5542.6,3120.2,10249.,1463.9,4802.0,736.14,2116.5,2586.9,0.0000,-4705.6,-7494.1,-427.15,-3378.8,-3301.8,-14651.,-1732.3,-1561.1,-5423.9,-3066.6,-5975.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
219.0000000000,36217.,2494.2,4417.5,6094.2,5554.5,3123.5,10261.,1459.8,4799.9,734.72,2110.5,2585.7,0.0000,-4696.6,-7485.9,-426.19,-3377.4,-3298.2,-14647.,-1732.2,-1557.7,-5423.0,-3066.5,-5973.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
220.0000000000,36231.,2438.7,4354.2,6030.7,5548.1,3122.1,10213.,1454.6,4791.1,733.06,2106.7,2567.4,0.0000,-4687.6,-7478.1,-425.25,-3375.9,-3294.6,-14643.,-1732.0,-1554.5,-5422.6,-3066.3,-5971.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
221.0000000000,36231.,2417.3,4239.3,6014.9,5549.0,3118.5,10155.,1454.7,4774.7,730.06,2090.9,2547.7,0.0000,-4679.1,-7470.4,-424.36,-3374.5,-3291.2,-14639.,-1731.9,-1551.6,-5421.9,-3066.0,-5969.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
222.0000000000,36219.,2430.6,4194.9,5980.5,5537.9,3118.1,10099.,1454.8,4754.1,728.29,2080.4,2543.5,0.0000,-4671.2,-7462.8,-423.49,-3373.0,-3287.9,-14635.,-1731.8,-1549.0,-5421.0,-3065.9,-5967.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
223.0000000000,36172.,2401.6,4175.2,5966.4,5470.1,3126.9,10096.,1457.0,4682.5,723.60,2077.0,2522.1,0.0000,-4663.4,-7456.0,-422.65,-3371.8,-3284.6,-14632.,-1731.9,-1546.4,-5420.4,-3065.7,-5966.0,1250.8,559.06,428.26,401.94,779.17,268.50,962.42,278.11,425.17,126.91,182.39,219.70,0.0000,-1.5246,-1.5944,-0.20249,-1.3357,-1.2814,-5.1542,-3.9985,-0.40497,-3.6005,-0.48321,-4.8867
224.0000000000,36165.,2374.4,4156.9,5968.9,5436.7,3132.0,10055.,1457.3,4686.1,717.06,2056.6,2500.2,0.0000,-4706.7,-7476.6,-426.10,-3370.8,-3309.7,-14629.,-1732.8,-1573.2,-5431.7,-3068.1,-5972.5,6864.2,3068.1,2350.3,2205.8,4276.1,1473.5,5281.7,1526.3,2333.3,696.47,1001.0,1205.7,0.0000,-8.3795,-8.7551,-1.1112,-7.3378,-7.0429,-28.276,-21.944,-2.2225,-19.759,-2.6520,-26.821
225.0000000000,36166.,2313.4,4085.0,5923.2,5422.8,3069.3,9948.9,1455.0,4672.9,713.47,2051.2,2496.0,0.0000,-4676.0,-7472.3,-424.97,-3369.7,-3289.1,-14624.,-1732.5,-1557.6,-5423.2,-3066.2,-5965.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
226.0000000000,36166.,2295.2,4067.7,5887.5,5374.5,3047.9,9911.0,1452.5,4618.4,708.19,2045.8,2468.4,0.0000,-4664.4,-7463.8,-423.42,-3368.8,-3283.7,-14620.,-1732.2,-1551.6,-5420.5,-3065.5,-5962.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
227.0000000000,36171.,2295.0,4028.8,5861.5,5318.6,3044.5,9861.5,1445.8,4617.1,706.30,2041.1,2443.0,0.0000,-4655.0,-7454.7,-422.03,-3367.8,-3279.7,-14616.,-1731.9,-1547.7,-5419.3,-3064.9,-5959.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
228.0000000000,36174.,2295.6,4028.6,5858.0,5273.0,3048.6,9833.5,1441.5,4590.6,705.92,2036.2,2434.7,0.0000,-4646.3,-7446.5,-420.83,-3366.6,-3276.1,-14612.,-1731.7,-1544.6,-5418.5,-3064.4,-5957.8,65.921,29.465,22.571,21.184,41.066,14.151,50.724,14.658,22.409,6.6887,9.6128,11.579,0.0000,-0.80148E-01,-0.83910E-01,-0.10672E-01,-0.70281E-01,-0.67252E-01,-0.27117,-0.21072,-0.21344E-01,-0.18972,-0.25458E-01,-0.25766
229.0000000000,35805.,2294.0,4022.4,5823.6,5244.5,3048.5,9810.0,1431.0,4571.8,702.96,2020.9,2425.4,0.0000,-4638.2,-7438.9,-419.78,-3365.5,-3272.8,-14608.,-1731.6,-1541.8,-5417.5,-3064.0,-5955.8,0.84258,0.37662,0.28850,0.27076,0.52489,0.18087,0.64834,0.18735,0.28642,0.85492E-01,0.12287,0.14800,0.0000,-0.10233E-02,-0.10718E-02,-0.13641E-03,-0.89778E-03,-0.85849E-03,-0.34647E-02,-0.26932E-02,-0.27281E-03,-0.24249E-02,-0.32534E-03,-0.32936E-02
230.0000000000,35531.,2274.3,3993.8,5775.9,5201.4,3009.2,9743.9,1430.0,4526.3,702.26,2010.3,2413.1,0.0000,-4630.4,-7431.8,-418.83,-3364.4,-3269.7,-14604.,-1731.4,-1539.2,-5416.7,-3063.5,-5953.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
231.0000000000,35439.,2258.4,3942.5,5722.0,5208.3,3009.3,9684.1,1423.2,4526.0,702.56,2014.2,2390.8,0.0000,-4622.9,-7424.9,-417.93,-3363.4,-3266.6,-14599.,-1731.3,-1536.8,-5415.9,-3063.2,-5952.1,103.13,46.096,35.311,33.140,64.244,22.138,79.353,22.931,35.056,10.464,15.038,18.114,0.0000,-0.12500,-0.13103,-0.16695E-01,-0.10976,-0.10481,-0.42377,-0.32960,-0.33391E-01,-0.29676,-0.39810E-01,-0.40317
232.0000000000,35444.,2262.0,3933.4,5660.4,5209.1,3001.2,9637.4,1414.1,4503.8,701.55,2015.0,2390.0,0.0000,-4615.6,-7418.1,-417.10,-3362.3,-3263.5,-14593.,-1731.2,-1534.6,-5415.2,-3063.0,-5950.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
233.0000000000,35333.,2224.0,3927.7,5636.2,5178.8,2988.8,9611.6,1395.1,4473.5,697.62,2014.0,2383.2,0.0000,-4608.3,-7411.7,-416.30,-3361.0,-3260.4,-14588.,-1731.1,-1532.4,-5414.5,-3062.9,-5948.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
234.0000000000,35280.,2231.2,3897.1,5634.3,5176.7,2935.8,9568.8,1382.1,4465.8,695.87,2014.2,2377.4,0.0000,-4651.5,-7432.3,-419.80,-3360.1,-3285.7,-14583.,-1731.6,-1559.2,-5425.4,-3065.5,-5954.8,4292.0,1918.5,1469.6,1379.3,2673.8,921.36,3302.6,954.37,1459.0,435.49,625.88,753.90,0.0000,-5.2000,-5.4502,-0.69484,-4.5683,-4.3582,-17.619,-13.715,-1.3897,-12.349,-1.6564,-16.783
235.0000000000,34773.,2189.4,3887.8,5629.4,5141.8,2912.9,9571.9,1375.8,4436.3,696.35,2006.1,2377.8,0.0000,-4620.8,-7428.8,-418.74,-3358.9,-3265.4,-14578.,-1731.4,-1544.1,-5416.8,-3063.8,-5947.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
236.0000000000,34596.,2173.5,3899.4,5630.0,5131.5,2931.4,9573.3,1365.4,4441.2,696.58,2005.7,2374.9,0.0000,-4659.7,-7448.1,-421.51,-3357.8,-3288.5,-14573.,-1746.7,-1567.7,-5428.8,-3065.8,-5957.1,0.11381E+06,50870.,38968.,36572.,70897.,24431.,87571.,25306.,38687.,11547.,16596.,19990.,0.0000,-137.95,-144.56,-18.424,-121.15,-115.53,-466.89,-363.66,-36.849,-327.41,-43.916,-445.10
237.0000000000,34561.,2143.5,3900.8,5604.5,5127.7,2939.9,9485.0,1363.3,4437.1,685.67,2008.0,2359.9,0.0000,-4677.7,-7469.2,-424.13,-3356.9,-3295.8,-14568.,-1743.2,-1580.3,-5432.5,-3066.6,-5959.8,2554.3,1141.7,874.58,820.83,1591.2,548.32,1965.4,567.96,868.28,259.17,372.47,448.66,0.0000,-3.1007,-3.2473,-0.41351,-2.7211,-2.5957,-10.476,-8.1617,-0.82703,-7.3483,-0.98566,-9.9908
238.0000000000,34427.,2128.9,3893.1,5552.7,5124.4,2948.3,9465.4,1360.8,4422.5,682.63,1993.0,2341.2,0.0000,-4691.9,-7488.6,-426.18,-3356.0,-3301.3,-14562.,-1742.1,-1589.7,-5433.4,-3067.0,-5960.0,16440.,7348.4,5629.1,5283.1,10241.,3529.2,12650.,3655.6,5588.5,1668.1,2397.4,2887.7,0.0000,-19.985,-20.919,-2.6615,-17.524,-16.722,-67.408,-52.530,-5.3230,-47.294,-6.3440,-64.311
239.0000000000,34369.,2121.7,3899.3,5540.7,5063.1,2950.8,9442.1,1362.0,4414.7,675.82,1984.5,2338.7,0.0000,-4704.4,-7505.9,-427.75,-3355.2,-3306.2,-14557.,-1759.0,-1597.5,-5437.1,-3067.2,-5963.9,0.14698E+06,65698.,50326.,47233.,91563.,31552.,0.11310E+06,32682.,49964.,14914.,21433.,25818.,0.0000,-178.91,-187.19,-23.795,-156.76,-149.63,-602.50,-469.70,-47.590,-422.82,-56.718,-575.06
240.0000000000,34234.,2122.3,3899.4,5516.5,4461.7,2976.2,9472.8,1364.8,4401.4,676.24,1973.0,2343.7,0.0000,-4715.3,-7521.4,-429.00,-3354.7,-3311.9,-14553.,-1768.0,-1604.5,-5441.7,-3067.4,-5968.7,0.11947E+06,53402.,40908.,38393.,74427.,25647.,91931.,26566.,40613.,12122.,17422.,20986.,0.0000,-145.64,-152.31,-19.342,-127.52,-121.84,-489.77,-381.88,-38.683,-343.72,-46.104,-467.64
241.0000000000,34211.,2195.5,3931.3,5510.5,4349.4,2980.6,9564.0,1389.3,4356.3,695.03,1992.2,2348.0,0.0000,-4679.5,-7511.3,-425.79,-3354.7,-3290.4,-14551.,-1758.3,-1580.4,-5431.8,-3067.3,-5960.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
242.0000000000,33990.,2237.6,3920.8,5483.9,4323.9,2951.4,9544.6,1388.8,4345.9,692.36,1990.3,2369.3,0.0000,-4665.1,-7499.3,-422.77,-3354.6,-3284.0,-14550.,-1750.6,-1569.8,-5429.8,-3068.4,-5954.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
243.0000000000,32806.,2203.6,3878.1,5462.7,4170.3,2931.3,9412.0,1371.2,4346.1,682.06,1984.2,2367.4,0.0000,-4652.5,-7484.3,-420.39,-3354.2,-3278.6,-14546.,-1744.9,-1562.6,-5427.3,-3070.2,-5950.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
244.0000000000,32784.,2152.6,3856.6,5408.3,4141.5,2917.2,9347.4,1375.4,4334.4,679.55,1977.2,2362.9,0.0000,-4640.5,-7469.6,-418.61,-3353.0,-3273.8,-14541.,-1740.9,-1556.8,-5424.3,-3070.6,-5945.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
245.0000000000,32717.,2120.2,3853.8,5387.5,4126.0,2871.1,9312.8,1376.1,4329.2,678.09,1984.1,2346.7,0.0000,-4629.3,-7458.2,-417.23,-3351.0,-3269.5,-14537.,-1738.0,-1551.9,-5421.9,-3072.0,-5942.2,61.720,27.587,21.133,19.834,38.449,13.249,47.491,13.724,20.980,6.2624,9.0001,10.841,0.0000,-0.74893E-01,-0.78467E-01,-0.99918E-02,-0.65678E-01,-0.62527E-01,-0.25302,-0.19776,-0.19984E-01,-0.17778,-0.23870E-01,-0.24210
246.0000000000,32602.,2087.3,3813.0,5394.7,4117.2,2879.8,9279.2,1365.5,4311.0,670.54,1993.1,2330.3,0.0000,-4668.9,-7474.2,-420.35,-3349.4,-3294.0,-14534.,-1743.1,-1577.2,-5433.0,-3076.8,-5948.7,51626.,23076.,17677.,16590.,32161.,11082.,39725.,11479.,17549.,5238.3,7528.3,9068.2,0.0000,-62.703,-65.655,-8.3578,-54.981,-52.358,-211.55,-165.42,-16.716,-148.70,-19.964,-202.54
247.0000000000,32476.,2062.5,3796.2,5387.1,4001.8,2862.9,9246.9,1363.1,4292.7,663.68,1969.0,2314.6,0.0000,-4636.4,-7466.2,-419.04,-3347.8,-3272.7,-14529.,-1739.9,-1559.7,-5423.6,-3076.3,-5941.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
248.0000000000,32464.,2010.1,3766.8,5322.7,3895.3,2870.1,9273.8,1364.9,4298.2,657.95,1938.8,2307.9,0.0000,-4673.9,-7480.8,-421.67,-3346.4,-3295.2,-14526.,-1743.0,-1581.8,-5432.3,-3078.2,-5947.3,40350.,18036.,13816.,12967.,25136.,8661.9,31048.,8972.2,13716.,4094.1,5884.0,7087.6,0.0000,-49.002,-51.318,-6.5323,-42.969,-40.887,-165.22,-129.29,-13.065,-116.21,-15.599,-158.33
249.0000000000,32385.,1986.3,3765.1,5291.6,3889.7,2870.6,9293.6,1355.5,4303.1,658.46,1914.4,2306.4,0.0000,-4690.2,-7498.2,-424.20,-3345.1,-3301.8,-14523.,-1743.3,-1592.8,-5434.4,-3078.4,-5948.6,24550.,10973.,8405.9,7889.2,15294.,5270.1,18890.,5458.9,8345.3,2491.0,3579.9,4312.2,0.0000,-29.851,-31.246,-3.9744,-26.160,-24.898,-100.49,-78.661,-7.9488,-70.705,-9.4898,-96.343
250.0000000000,32345.,1968.3,3759.9,5227.0,3865.2,2854.9,9298.5,1355.1,4290.3,659.89,1891.3,2302.0,0.0000,-4652.3,-7487.8,-421.93,-3343.7,-3278.1,-14519.,-1740.0,-1570.8,-5422.7,-3076.0,-5939.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
251.0000000000,32222.,1914.7,3753.9,5216.5,3845.0,2852.1,9216.4,1345.1,4283.9,659.63,1883.1,2293.7,0.0000,-4636.5,-7473.0,-419.51,-3342.1,-3271.1,-14516.,-1737.5,-1561.4,-5418.4,-3074.7,-5935.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
252.0000000000,32077.,1875.9,3765.6,5206.1,3822.6,2842.9,9187.3,1338.8,4220.3,659.36,1876.0,2297.6,0.0000,-4675.1,-7485.7,-421.80,-3341.0,-3294.8,-14514.,-1740.1,-1584.5,-5428.2,-3076.2,-5941.1,32719.,14625.,11203.,10514.,20383.,7023.8,25176.,7275.4,11122.,3319.9,4771.2,5747.2,0.0000,-39.730,-41.625,-5.2970,-34.830,-33.109,-133.83,-104.83,-10.594,-94.226,-12.642,-128.45
253.0000000000,31891.,1809.8,3767.3,5151.7,3768.4,2834.6,9098.3,1339.6,4203.9,658.27,1851.4,2289.1,0.0000,-4692.2,-7502.1,-424.16,-3340.3,-3301.6,-14511.,-1738.5,-1595.4,-5430.6,-3076.1,-5942.3,5496.2,2456.7,1881.9,1766.2,3423.9,1179.9,4229.1,1222.1,1868.3,557.67,801.47,965.41,0.0000,-6.6839,-6.9978,-0.88978,-5.8550,-5.5685,-22.476,-17.610,-1.7796,-15.829,-2.1239,-21.581
254.0000000000,31801.,1816.2,3709.6,5153.9,3720.2,2838.0,9047.3,1340.5,4163.4,656.36,1821.2,2281.1,0.0000,-4704.8,-7517.6,-426.04,-3339.5,-3306.4,-14509.,-1738.7,-1603.0,-5431.2,-3075.6,-5942.1,16232.,7255.2,5557.7,5216.1,10112.,3484.4,12490.,3609.2,5517.6,1646.9,2367.0,2851.1,0.0000,-19.765,-20.683,-2.6278,-17.301,-16.461,-66.364,-52.012,-5.2555,-46.748,-6.2730,-63.742
255.0000000000,30795.,1809.1,3672.3,5150.0,3715.1,2819.1,8994.7,1338.3,4077.5,656.30,1801.1,2280.0,0.0000,-4664.5,-7504.0,-423.22,-3338.4,-3282.0,-14506.,-1736.7,-1579.0,-5419.6,-3072.9,-5933.0,159.47,71.279,54.602,51.246,99.342,34.233,122.71,35.459,54.208,16.181,23.254,28.011,0.0000,-0.19392,-0.20311,-0.25817E-01,-0.16979,-0.16141,-0.65180,-0.51099,-0.51633E-01,-0.45927,-0.61620E-01,-0.62630
256.0000000000,30493.,1799.9,3620.3,5148.8,3711.8,2810.6,8958.9,1337.8,4053.5,654.98,1800.8,2277.2,0.0000,-4646.6,-7486.7,-420.42,-3337.3,-3274.7,-14503.,-1735.1,-1568.5,-5415.5,-3072.5,-5928.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
257.0000000000,30475.,1798.3,3595.6,5124.9,3694.9,2818.8,8902.7,1330.5,4007.1,650.11,1780.7,2256.4,0.0000,-4632.5,-7470.6,-418.17,-3336.1,-3269.4,-14500.,-1733.9,-1561.2,-5413.5,-3072.4,-5926.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
258.0000000000,30471.,1774.8,3558.7,5033.1,3624.3,2815.8,8863.0,1330.1,3991.5,648.73,1766.5,2257.5,0.0000,-4619.9,-7456.4,-416.40,-3334.7,-3264.9,-14496.,-1733.0,-1555.2,-5412.0,-3072.3,-5924.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
259.0000000000,30413.,1752.2,3528.3,4999.0,3520.4,2812.7,8850.9,1329.6,3998.1,634.37,1768.2,2255.1,0.0000,-4608.6,-7443.2,-414.96,-3333.3,-3260.8,-14493.,-1732.4,-1550.5,-5410.8,-3072.4,-5922.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
260.0000000000,30354.,1726.9,3517.5,5000.8,3494.8,2806.9,8789.9,1327.0,4008.7,627.28,1758.9,2245.3,0.0000,-4649.0,-7458.0,-418.01,-3332.5,-3285.5,-14491.,-1735.7,-1575.7,-5422.1,-3075.3,-5929.5,27762.,12409.,9505.6,8921.4,17294.,5959.6,21362.,6173.0,9437.1,2816.9,4048.3,4876.4,0.0000,-33.618,-35.272,-4.4944,-29.497,-27.977,-113.34,-88.937,-8.9888,-79.940,-10.724,-109.08
261.0000000000,30294.,1718.9,3490.3,4995.1,3465.3,2817.0,8798.3,1324.4,4013.5,627.90,1753.0,2208.7,0.0000,-4666.7,-7476.2,-420.90,-3332.1,-3292.9,-14489.,-1741.9,-1588.0,-5427.0,-3076.9,-5932.9,54245.,24247.,18574.,17432.,33792.,11645.,41740.,12062.,18440.,5504.0,7910.2,9528.3,0.0000,-65.780,-68.968,-8.7818,-57.678,-54.730,-221.41,-173.78,-17.564,-156.19,-20.956,-213.16
262.0000000000,30246.,1706.5,3489.1,4995.5,3446.4,2809.8,8807.9,1322.6,4012.7,630.94,1740.3,2191.4,0.0000,-4680.5,-7493.7,-423.13,-3331.7,-3298.0,-14487.,-1740.8,-1596.7,-5429.4,-3077.6,-5934.0,12709.,5680.9,4351.7,4084.2,7917.4,2728.3,9779.5,2826.0,4320.3,1289.6,1853.3,2232.4,0.0000,-15.432,-16.171,-2.0575,-13.522,-12.834,-51.865,-40.715,-4.1151,-36.594,-4.9097,-49.947
263.0000000000,30225.,1693.4,3492.8,4992.5,3439.9,2811.6,8808.4,1314.8,4002.1,630.33,1719.9,2170.4,0.0000,-4693.0,-7509.0,-424.82,-3331.2,-3302.2,-14485.,-1782.3,-1603.8,-5439.0,-3077.5,-5945.0,0.32489E+06,0.14522E+06,0.11124E+06,0.10440E+06,0.20239E+06,69742.,0.24999E+06,72241.,0.11044E+06,32965.,47376.,57067.,0.0000,-395.00,-413.67,-52.596,-345.84,-328.34,-1325.7,-1041.1,-105.19,-935.44,-125.50,-1277.0
264.0000000000,30226.,1852.7,3607.5,4989.7,3475.1,2930.6,9007.1,1351.6,3948.5,673.19,1768.8,2209.7,0.0000,-4714.1,-7529.8,-426.25,-3333.2,-3313.8,-14490.,-1805.6,-1610.0,-5453.0,-3081.8,-5958.7,0.26417E+06,0.11808E+06,90450.,84890.,0.16456E+06,56708.,0.20327E+06,58739.,89798.,26804.,38521.,46401.,0.0000,-322.95,-337.26,-42.766,-282.00,-268.67,-1080.4,-848.35,-85.532,-761.68,-102.39,-1040.2
265.0000000000,30207.,2007.7,3679.4,4987.3,3521.2,2893.5,9039.6,1370.1,3945.7,700.60,1846.5,2297.6,0.0000,-4689.7,-7526.2,-423.35,-3339.2,-3294.2,-14499.,-1786.1,-1584.9,-5454.5,-3090.9,-5954.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
266.0000000000,30197.,2014.5,3699.7,4980.7,3574.5,2888.3,8877.0,1379.6,3992.0,707.37,1969.9,2300.1,0.0000,-4677.9,-7520.6,-420.82,-3340.6,-3287.8,-14504.,-1771.0,-1575.0,-5453.0,-3108.7,-5950.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
267.0000000000,30255.,1885.1,3627.0,4943.0,3505.0,2878.5,8943.9,1365.6,3994.8,687.60,1910.0,2236.4,0.0000,-4670.5,-7507.2,-418.93,-3338.4,-3281.4,-14507.,-1759.6,-1568.3,-5446.1,-3117.8,-5945.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
268.0000000000,30120.,1842.3,3650.2,4948.6,3565.2,2857.5,9017.9,1342.2,3999.8,690.26,1805.9,2217.1,0.0000,-4662.1,-7489.1,-417.45,-3336.1,-3275.2,-14508.,-1751.5,-1562.6,-5440.9,-3116.4,-5940.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
269.0000000000,29609.,1729.6,3628.7,4920.6,3684.8,2832.3,8867.0,1334.1,3997.1,690.40,1768.7,2220.8,0.0000,-4652.0,-7473.7,-416.26,-3334.2,-3270.2,-14509.,-1745.8,-1557.6,-5436.6,-3111.9,-5937.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
270.0000000000,29582.,1654.8,3615.1,4888.1,3597.6,2835.2,8795.9,1329.3,3955.9,687.75,1802.2,2222.8,0.0000,-4640.5,-7461.8,-415.22,-3333.0,-3265.8,-14508.,-1741.9,-1553.2,-5433.3,-3113.2,-5935.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
271.0000000000,29573.,1634.7,3667.4,4881.8,3566.5,2856.2,8836.9,1316.4,3968.8,687.23,1762.6,2220.3,0.0000,-4631.7,-7452.2,-414.27,-3332.0,-3261.6,-14508.,-1739.2,-1550.8,-5431.8,-3112.2,-5934.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
272.0000000000,29532.,1622.6,3647.8,4890.9,3648.0,2907.1,8846.0,1304.4,3950.1,682.59,1748.0,2198.2,0.0000,-4675.0,-7467.6,-417.63,-3334.5,-3286.4,-14510.,-1743.4,-1577.4,-5445.1,-3111.1,-5941.5,44135.,19728.,15112.,14183.,27494.,9474.4,33961.,9813.8,15003.,4478.2,6435.9,7752.4,0.0000,-53.594,-56.144,-7.1451,-46.967,-44.552,-180.26,-142.17,-14.290,-127.52,-17.124,-174.25
273.0000000000,29534.,1642.0,3630.1,4889.2,3572.0,2907.6,8789.6,1291.3,3910.7,680.55,1700.6,2176.6,0.0000,-4643.1,-7461.3,-416.48,-3335.6,-3265.5,-14508.,-1740.6,-1560.6,-5436.5,-3106.2,-5934.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
274.0000000000,29476.,1576.8,3631.8,4866.1,3555.0,2890.8,8739.6,1290.7,3903.7,672.09,1690.9,2180.5,0.0000,-4630.1,-7452.9,-414.91,-3338.0,-3261.2,-14506.,-1738.5,-1553.8,-5433.3,-3103.8,-5931.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
275.0000000000,29470.,1563.5,3617.7,4811.7,3544.2,2872.9,8691.8,1294.6,3910.8,675.95,1696.7,2166.0,0.0000,-4619.3,-7443.5,-413.54,-3340.2,-3258.0,-14504.,-1736.9,-1549.2,-5431.0,-3103.2,-5928.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
276.0000000000,29445.,1613.3,3605.1,4775.8,3551.5,2865.3,8672.7,1301.5,3877.9,672.88,1699.1,2140.0,0.0000,-4609.7,-7435.0,-412.39,-3342.0,-3254.9,-14502.,-1735.7,-1545.3,-5429.1,-3103.3,-5926.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
277.0000000000,29393.,1621.7,3564.6,4785.6,3547.7,2885.6,8670.7,1298.4,3883.1,673.35,1685.5,2133.5,0.0000,-4600.9,-7427.0,-411.41,-3343.1,-3251.8,-14502.,-1734.9,-1542.1,-5427.7,-3102.3,-5924.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
278.0000000000,29324.,1607.6,3517.6,4736.7,3520.5,2888.2,8585.4,1287.4,3902.3,671.69,1689.5,2123.2,0.0000,-4592.7,-7417.8,-410.54,-3344.1,-3248.9,-14500.,-1734.3,-1539.2,-5426.1,-3100.8,-5922.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
279.0000000000,29279.,1596.9,3523.7,4715.2,3434.8,2862.6,8587.0,1288.7,3889.7,671.83,1680.7,2097.0,0.0000,-4583.7,-7409.1,-409.77,-3344.6,-3245.8,-14500.,-1733.9,-1536.0,-5424.8,-3099.8,-5920.3,439.44,196.42,150.47,141.22,273.75,94.334,338.14,97.714,149.38,44.588,64.081,77.189,0.0000,-0.52968,-0.55690,-0.71142E-01,-0.46619,-0.44064,-1.7922,-1.4136,-0.14228,-1.2684,-0.17027,-1.7351
280.0000000000,28661.,1562.6,3526.8,4723.9,3399.3,2792.7,8544.5,1294.7,3892.9,662.45,1681.3,2089.8,0.0000,-4574.8,-7402.0,-409.09,-3344.5,-3242.8,-14499.,-1733.5,-1533.3,-5422.4,-3099.2,-5918.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
281.0000000000,28325.,1507.8,3507.8,4701.3,3391.2,2768.5,8538.3,1302.8,3882.5,657.47,1691.8,2091.1,0.0000,-4566.2,-7395.7,-408.44,-3344.3,-3239.8,-14498.,-1733.3,-1531.0,-5421.1,-3098.8,-5917.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
282.0000000000,27982.,1502.1,3517.3,4679.4,3339.5,2754.8,8479.1,1301.7,3876.8,661.52,1668.7,2093.3,0.0000,-4557.9,-7387.8,-407.83,-3343.1,-3235.6,-14496.,-1733.1,-1528.8,-5420.4,-3098.1,-5916.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
283.0000000000,27870.,1438.6,3534.1,4676.3,3311.9,2762.8,8447.1,1296.8,3850.6,658.43,1647.1,2096.9,0.0000,-4549.7,-7380.9,-407.23,-3342.0,-3231.8,-14494.,-1732.9,-1526.8,-5419.8,-3096.6,-5915.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
284.0000000000,27241.,1412.3,3503.8,4674.8,3247.8,2752.0,8344.3,1285.5,3859.8,658.37,1637.4,2084.1,0.0000,-4541.7,-7374.4,-406.65,-3341.1,-3228.2,-14492.,-1732.8,-1524.7,-5419.5,-3095.3,-5914.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
285.0000000000,27124.,1432.0,3504.1,4651.3,3188.9,2719.8,8328.7,1275.5,3859.2,660.17,1624.6,2073.6,0.0000,-4534.0,-7368.4,-406.08,-3340.1,-3224.7,-14490.,-1732.7,-1522.5,-5419.2,-3093.9,-5914.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
286.0000000000,27095.,1394.2,3436.7,4665.8,3095.3,2749.7,8382.1,1264.6,3866.5,665.49,1618.8,2066.9,0.0000,-4526.6,-7362.1,-405.53,-3339.1,-3221.3,-14490.,-1732.7,-1520.6,-5418.6,-3092.7,-5913.5,1181.3,528.02,404.48,379.62,735.90,253.59,908.98,262.67,401.56,119.86,172.26,207.50,0.0000,-1.4137,-1.4922,-0.19124,-1.2502,-1.1766,-4.8119,-3.7952,-0.38249,-3.4073,-0.45848,-4.6649
287.0000000000,27010.,1397.3,3395.9,4690.8,3017.4,2784.1,8395.1,1246.5,3863.1,670.34,1593.8,2053.7,0.0000,-4569.2,-7380.4,-409.23,-3338.3,-3246.3,-14492.,-1738.0,-1547.6,-5430.7,-3094.4,-5922.3,39533.,17670.,13536.,12704.,24627.,8486.4,30419.,8790.4,13438.,4011.2,5764.8,6944.0,0.0000,-47.383,-49.970,-6.4000,-41.881,-39.448,-161.00,-126.99,-12.800,-114.02,-15.348,-156.12
288.0000000000,26903.,1367.7,3381.1,4685.5,2980.1,2772.4,8426.9,1242.8,3866.2,658.70,1579.7,2043.4,0.0000,-4588.7,-7401.0,-412.64,-3337.5,-3254.1,-14492.,-1746.5,-1562.9,-5436.1,-3095.2,-5927.5,72001.,32183.,24653.,23138.,44853.,15456.,55402.,16010.,24475.,7305.5,10499.,12647.,0.0000,-86.441,-91.093,-11.656,-76.338,-71.953,-293.17,-231.26,-23.312,-207.64,-27.960,-284.34
289.0000000000,26902.,1347.4,3347.2,4674.8,2907.6,2768.0,8382.2,1245.5,3789.5,648.74,1577.1,2023.6,0.0000,-4603.7,-7420.8,-415.27,-3336.8,-3259.8,-14491.,-1772.8,-1574.2,-5443.8,-3095.5,-5937.0,0.21906E+06,97915.,75005.,70395.,0.13646E+06,47025.,0.16856E+06,48709.,74464.,22227.,31944.,38478.,0.0000,-263.41,-277.41,-35.463,-232.40,-219.19,-891.79,-703.65,-70.927,-631.70,-85.079,-865.18
290.0000000000,26901.,1397.3,3336.8,4720.7,2924.2,2772.4,8422.3,1254.4,3768.7,661.18,1570.3,2025.0,0.0000,-4619.6,-7439.1,-417.31,-3337.0,-3268.0,-14492.,-1763.5,-1583.7,-5446.9,-3096.6,-5941.0,5396.8,2412.3,1847.9,1734.3,3362.0,1158.5,4152.7,1200.0,1834.5,547.59,786.98,947.96,0.0000,-6.5087,-6.8459,-0.87370,-5.7345,-5.4199,-21.989,-17.343,-1.7474,-15.570,-2.0982,-21.331
291.0000000000,26664.,1451.3,3329.9,4737.8,2901.8,2711.4,8431.1,1269.6,3711.3,664.70,1571.4,2022.0,0.0000,-4585.5,-7434.5,-414.66,-3336.7,-3245.4,-14495.,-1755.1,-1562.2,-5436.4,-3096.4,-5932.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
292.0000000000,26209.,1434.5,3285.9,4761.8,2885.0,2685.7,8323.9,1259.1,3733.2,654.11,1567.6,2011.7,0.0000,-4572.1,-7420.2,-412.02,-3338.3,-3238.4,-14494.,-1748.9,-1553.8,-5432.4,-3097.3,-5927.0,1034.7,462.47,354.27,332.49,644.55,222.11,796.14,230.06,351.71,104.98,150.88,181.74,0.0000,-1.2465,-1.3115,-0.16750,-1.0978,-1.0363,-4.2171,-3.3280,-0.33500,-2.9870,-0.40277,-4.0920
293.0000000000,26081.,1403.2,3260.3,4740.3,2820.1,2661.8,8232.2,1261.9,3725.8,647.38,1570.0,1995.8,0.0000,-4560.1,-7405.4,-409.94,-3338.7,-3233.2,-14489.,-1744.2,-1548.5,-5428.8,-3097.2,-5923.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
294.0000000000,26055.,1367.0,3267.1,4734.8,2797.6,2655.1,8236.9,1262.2,3701.5,641.16,1576.5,1970.0,0.0000,-4549.3,-7394.0,-408.36,-3338.5,-3229.0,-14485.,-1740.9,-1544.0,-5425.8,-3098.6,-5919.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
295.0000000000,26063.,1394.5,3275.4,4718.9,2792.2,2660.9,8243.5,1261.1,3695.4,639.25,1570.6,1944.2,0.0000,-4539.0,-7383.3,-407.12,-3337.9,-3225.3,-14481.,-1738.6,-1540.1,-5423.9,-3100.3,-5916.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
296.0000000000,26045.,1360.3,3259.9,4647.6,2707.0,2718.9,8235.3,1266.4,3688.1,622.89,1575.6,1933.0,0.0000,-4529.5,-7374.0,-406.07,-3337.1,-3221.4,-14478.,-1737.0,-1536.6,-5422.3,-3101.9,-5913.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
297.0000000000,26059.,1320.2,3275.7,4583.4,2711.3,2747.8,8143.9,1263.4,3622.3,618.16,1560.8,1928.1,0.0000,-4521.2,-7366.2,-405.14,-3336.3,-3217.5,-14471.,-1735.8,-1533.4,-5421.4,-3102.2,-5911.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
298.0000000000,25495.,1312.2,3287.3,4551.3,2686.0,2735.4,8111.3,1255.9,3532.0,616.20,1535.5,1907.6,0.0000,-4512.9,-7359.8,-404.31,-3334.4,-3213.9,-14464.,-1735.0,-1530.3,-5420.0,-3101.3,-5909.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
299.0000000000,25007.,1289.9,3307.2,4486.7,2665.1,2725.7,8064.2,1263.2,3531.7,615.56,1518.1,1890.6,0.0000,-4505.3,-7353.7,-403.56,-3332.3,-3210.9,-14458.,-1734.4,-1527.3,-5418.5,-3100.7,-5907.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
300.0000000000,24219.,1277.7,3314.3,4430.0,2654.7,2703.0,8028.2,1271.1,3548.4,619.82,1514.1,1871.5,0.0000,-4497.8,-7347.8,-402.86,-3330.2,-3208.1,-14452.,-1733.9,-1524.7,-5417.0,-3099.6,-5906.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
301.0000000000,23497.,1331.9,3300.5,4410.9,2658.4,2677.7,7991.4,1267.8,3507.7,625.74,1511.1,1842.3,0.0000,-4490.8,-7341.9,-402.21,-3328.2,-3205.4,-14447.,-1733.6,-1522.4,-5415.9,-3098.5,-5904.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
302.0000000000,22614.,1300.5,3269.4,4397.4,2628.6,2676.1,7941.8,1254.5,3472.2,619.27,1493.4,1838.6,0.0000,-4484.1,-7334.7,-401.58,-3326.4,-3202.6,-14443.,-1733.3,-1520.2,-5414.2,-3097.8,-5902.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
303.0000000000,22085.,1285.0,3265.8,4387.8,2608.5,2659.7,7907.2,1240.8,3420.4,613.73,1477.8,1813.1,0.0000,-4477.6,-7326.9,-400.96,-3324.7,-3199.5,-14439.,-1733.1,-1518.2,-5412.5,-3097.0,-5901.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
304.0000000000,21169.,1299.5,3289.9,4358.7,2542.6,2695.3,7883.9,1228.1,3363.5,590.36,1456.6,1784.2,0.0000,-4520.5,-7345.2,-404.58,-3323.5,-3224.5,-14436.,-1733.3,-1544.5,-5422.7,-3098.7,-5908.1,1822.6,814.67,624.06,585.70,1135.4,391.25,1402.4,405.27,619.56,184.93,265.78,320.14,0.0000,-2.1700,-2.2924,-0.29506,-1.9231,-1.8002,-7.4092,-5.8518,-0.59013,-5.2558,-0.70853,-7.2097
305.0000000000,20508.,1254.6,3316.0,4329.4,2531.5,2698.1,7857.6,1212.7,3330.5,582.57,1427.0,1764.1,0.0000,-4490.3,-7340.7,-403.67,-3322.2,-3203.7,-14433.,-1733.1,-1529.5,-5413.7,-3096.2,-5901.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
306.0000000000,20439.,1241.1,3343.3,4322.5,2520.8,2633.4,7844.3,1217.1,3362.3,584.65,1412.1,1765.2,0.0000,-4478.7,-7333.6,-402.31,-3320.8,-3198.1,-14430.,-1732.9,-1523.7,-5411.0,-3094.5,-5899.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
307.0000000000,20343.,1218.8,3328.8,4325.1,2504.2,2629.8,7846.9,1215.9,3355.2,581.73,1404.9,1757.8,0.0000,-4469.4,-7326.4,-401.10,-3319.0,-3194.0,-14429.,-1732.7,-1520.1,-5409.6,-3093.3,-5898.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
308.0000000000,20297.,1218.2,3306.5,4352.5,2498.8,2654.9,7801.3,1219.8,3356.1,584.22,1389.0,1748.4,0.0000,-4510.6,-7345.3,-404.42,-3317.6,-3218.8,-14428.,-1736.5,-1546.3,-5420.6,-3095.6,-5906.7,28299.,12649.,9689.7,9094.1,17629.,6074.9,21775.,6292.6,9619.8,2871.4,4126.7,4970.8,0.0000,-33.641,-35.559,-4.5814,-29.829,-27.874,-114.93,-90.788,-9.1628,-81.570,-10.998,-111.94
309.0000000000,20277.,1252.7,3274.1,4352.7,2491.8,2645.4,7755.8,1212.1,3383.2,581.49,1371.3,1728.9,0.0000,-4529.1,-7367.3,-407.61,-3316.5,-3226.6,-14427.,-1736.6,-1560.3,-5423.4,-3096.4,-5909.6,7881.6,3522.9,2698.7,2532.8,4909.9,1691.9,6064.7,1752.5,2679.2,799.71,1149.3,1384.4,0.0000,-9.3837,-9.9114,-1.2760,-8.3141,-7.7730,-32.001,-25.281,-2.5519,-22.716,-3.0634,-31.176
310.0000000000,20295.,1273.5,3252.7,4371.8,2459.7,2654.4,7743.2,1215.1,3369.4,580.74,1370.1,1737.9,0.0000,-4543.3,-7386.2,-410.12,-3315.6,-3232.3,-14425.,-1738.7,-1570.8,-5424.9,-3097.0,-5911.4,23784.,10631.,8143.7,7643.2,14817.,5105.7,18301.,5288.6,8085.0,2413.3,3468.3,4177.8,0.0000,-28.359,-29.935,-3.8505,-25.106,-23.481,-96.549,-76.275,-7.7009,-68.543,-9.2451,-94.080
311.0000000000,20283.,1302.7,3247.1,4300.7,2415.7,2644.1,7692.5,1213.1,3380.8,582.97,1351.3,1734.9,0.0000,-4555.7,-7403.5,-412.01,-3314.7,-3237.2,-14423.,-1739.7,-1579.3,-5425.7,-3097.3,-5912.9,19613.,8766.5,6715.3,6302.6,12218.,4210.2,15091.,4361.0,6666.9,1990.0,2860.0,3445.0,0.0000,-23.418,-24.706,-3.1751,-20.714,-19.379,-79.600,-62.886,-6.3502,-56.515,-7.6242,-77.579
312.0000000000,20281.,1271.4,3226.0,4256.5,2421.1,2613.7,7645.2,1199.5,3311.7,584.65,1326.7,1724.1,0.0000,-4516.5,-7392.2,-409.20,-3313.6,-3213.3,-14418.,-1737.7,-1557.3,-5414.0,-3094.8,-5905.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
313.0000000000,19714.,1236.6,3242.4,4236.5,2442.3,2556.3,7646.3,1182.4,3291.3,586.86,1324.7,1684.8,0.0000,-4550.3,-7402.8,-410.66,-3312.6,-3234.9,-14414.,-1739.3,-1577.3,-5421.9,-3096.4,-5910.9,22853.,10215.,7825.0,7344.0,14237.,4905.9,17585.,5081.6,7768.6,2318.8,3332.6,4014.2,0.0000,-27.285,-28.791,-3.6998,-24.129,-22.557,-92.723,-73.250,-7.3995,-65.841,-8.8847,-90.397
314.0000000000,19612.,1198.9,3284.2,4158.5,2485.8,2514.7,7639.1,1178.2,3221.5,580.52,1315.3,1676.0,0.0000,-4514.1,-7390.0,-408.12,-3311.2,-3212.5,-14409.,-1737.3,-1557.4,-5412.1,-3094.2,-5903.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
315.0000000000,19491.,1205.0,3272.9,4097.9,2467.9,2506.1,7631.0,1177.1,3190.6,573.06,1318.6,1674.3,0.0000,-4498.3,-7374.6,-405.62,-3309.8,-3206.0,-14405.,-1735.8,-1548.4,-5408.9,-3093.2,-5900.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
316.0000000000,18813.,1213.2,3269.0,4106.2,2431.8,2536.4,7507.0,1179.3,3191.2,563.14,1321.0,1652.7,0.0000,-4535.8,-7386.3,-407.84,-3308.7,-3229.7,-14402.,-1735.4,-1571.5,-5419.1,-3095.0,-5906.6,4693.6,2098.0,1607.1,1508.3,2923.9,1007.6,3611.6,1043.7,1595.5,476.24,684.44,824.44,0.0000,-5.5959,-5.9078,-0.75985,-4.9509,-4.6217,-19.035,-15.035,-1.5197,-13.518,-1.8246,-18.566
317.0000000000,18803.,1248.3,3231.0,4062.0,2402.9,2542.5,7446.8,1175.7,3193.6,556.39,1315.5,1638.8,0.0000,-4501.6,-7375.6,-405.93,-3307.4,-3208.4,-14397.,-1734.5,-1553.0,-5410.0,-3092.7,-5899.6,1138.2,508.75,389.72,365.76,709.05,244.33,875.81,253.09,386.91,115.49,165.98,199.93,0.0000,-1.3554,-1.4318,-0.18426,-1.1995,-1.1189,-4.6154,-3.6453,-0.36853,-3.2778,-0.44243,-4.5024
318.0000000000,18775.,1247.4,3230.7,3999.0,2404.1,2542.8,7442.0,1174.2,3144.1,556.51,1294.6,1623.4,0.0000,-4487.5,-7362.0,-403.86,-3306.0,-3202.4,-14393.,-1733.7,-1544.9,-5406.9,-3091.1,-5896.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
319.0000000000,18044.,1238.9,3234.0,3950.4,2380.5,2591.2,7422.4,1181.6,3094.0,547.09,1278.6,1603.2,0.0000,-4476.6,-7349.0,-402.15,-3304.5,-3197.9,-14390.,-1733.1,-1539.3,-5405.2,-3089.9,-5894.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
320.0000000000,17983.,1259.3,3253.3,3890.0,2357.1,2542.8,7277.5,1182.5,3116.8,545.15,1279.3,1584.7,0.0000,-4466.9,-7337.9,-400.76,-3303.0,-3193.9,-14387.,-1732.7,-1534.6,-5403.8,-3088.8,-5893.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
321.0000000000,17521.,1214.9,3266.6,3872.0,2354.1,2481.1,7228.0,1169.9,3107.4,540.14,1283.6,1579.3,0.0000,-4457.6,-7327.6,-399.60,-3301.9,-3190.5,-14383.,-1732.3,-1530.4,-5402.6,-3088.0,-5891.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
322.0000000000,17156.,1202.4,3254.6,3838.2,2342.1,2444.0,7132.9,1162.4,3075.5,539.27,1278.2,1563.5,0.0000,-4448.5,-7318.0,-398.60,-3300.7,-3187.0,-14380.,-1732.0,-1526.3,-5401.9,-3087.3,-5889.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
323.0000000000,17157.,1203.8,3247.1,3816.5,2342.5,2438.4,7034.7,1161.7,3065.9,540.40,1259.5,1547.9,0.0000,-4439.3,-7308.8,-397.72,-3299.3,-3183.4,-14377.,-1731.8,-1522.7,-5401.4,-3086.9,-5888.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
324.0000000000,17155.,1220.5,3245.1,3791.0,2332.5,2437.6,6956.1,1159.6,3070.4,538.80,1255.5,1528.2,0.0000,-4430.6,-7300.0,-396.92,-3297.4,-3179.9,-14373.,-1731.6,-1519.4,-5400.7,-3086.6,-5887.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
325.0000000000,17148.,1234.0,3242.3,3760.7,2308.8,2437.9,6909.0,1156.5,3074.0,539.22,1247.2,1516.7,0.0000,-4422.7,-7292.0,-396.19,-3295.7,-3176.6,-14370.,-1731.4,-1516.5,-5399.5,-3086.3,-5886.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
326.0000000000,17162.,1251.8,3247.0,3754.0,2271.8,2409.4,6871.4,1155.2,3059.8,541.04,1245.1,1495.0,0.0000,-4464.3,-7309.8,-399.72,-3294.3,-3201.5,-14367.,-1732.6,-1542.3,-5410.4,-3088.8,-5893.2,8980.8,4014.3,3075.0,2886.0,5594.7,1927.9,6910.5,1997.0,3052.9,911.24,1309.6,1577.5,0.0000,-10.611,-11.230,-1.4539,-9.4289,-8.7425,-36.364,-28.721,-2.9078,-25.849,-3.4885,-35.527
327.0000000000,16655.,1252.0,3257.2,3694.9,2248.8,2416.8,6806.3,1152.6,3056.4,542.56,1243.8,1477.2,0.0000,-4482.9,-7330.4,-402.99,-3293.0,-3209.3,-14364.,-1733.4,-1555.8,-5413.6,-3089.7,-5895.4,8660.3,3871.0,2965.3,2783.0,5395.0,1859.1,6663.8,1925.7,2943.9,878.71,1262.9,1521.2,0.0000,-10.248,-10.837,-1.4020,-9.0997,-8.4397,-35.058,-27.692,-2.8040,-24.925,-3.3642,-34.259
328.0000000000,16518.,1257.0,3258.2,3638.6,2165.0,2415.4,6760.7,1144.0,3062.7,542.85,1236.4,1469.2,0.0000,-4497.4,-7349.0,-405.53,-3291.9,-3214.9,-14361.,-1740.7,-1565.7,-5416.1,-3090.0,-5898.2,58339.,26077.,19975.,18748.,36343.,12524.,44890.,12972.,19831.,5919.4,8507.2,10247.,0.0000,-69.135,-73.059,-9.4446,-61.339,-56.902,-236.12,-186.52,-18.889,-167.90,-22.662,-230.78
329.0000000000,16517.,1249.5,3264.2,3639.3,2103.7,2421.4,6667.3,1132.7,3061.5,541.07,1227.8,1463.6,0.0000,-4509.8,-7364.6,-407.46,-3290.3,-3219.4,-14359.,-1744.6,-1574.0,-5418.3,-3090.1,-5900.9,46803.,20920.,16025.,15040.,29156.,10047.,36013.,10407.,15910.,4748.9,6825.0,8221.0,0.0000,-55.539,-58.657,-7.5770,-49.234,-45.682,-189.39,-149.62,-15.154,-134.69,-18.181,-185.15
330.0000000000,16518.,1232.7,3247.8,3636.9,2040.2,2412.4,6600.3,1120.2,3053.1,539.58,1216.5,1466.4,0.0000,-4471.0,-7352.4,-404.73,-3288.4,-3195.2,-14355.,-1741.2,-1551.6,-5407.2,-3087.4,-5893.3,1016.4,454.31,348.01,326.62,633.16,218.19,782.08,226.00,345.50,103.13,148.21,178.53,0.0000,-1.2046,-1.2732,-0.16454,-1.0680,-0.98978,-4.1120,-3.2487,-0.32909,-2.9248,-0.39475,-4.0207
331.0000000000,15956.,1225.1,3233.2,3636.4,2032.9,2410.5,6586.1,1117.9,3062.6,535.71,1208.2,1450.8,0.0000,-4454.4,-7337.0,-402.01,-3286.3,-3188.1,-14352.,-1738.3,-1542.1,-5403.0,-3085.9,-5889.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
332.0000000000,15871.,1222.8,3241.2,3611.8,2034.4,2406.1,6560.4,1114.0,3032.3,533.95,1204.6,1452.9,0.0000,-4441.5,-7322.2,-399.83,-3284.4,-3183.7,-14349.,-1736.0,-1535.6,-5400.3,-3084.6,-5886.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
333.0000000000,15824.,1229.2,3249.7,3581.6,2037.1,2404.7,6505.6,1114.2,3012.2,533.75,1182.5,1451.0,0.0000,-4430.9,-7308.6,-398.13,-3282.6,-3180.1,-14346.,-1734.4,-1530.3,-5398.4,-3083.9,-5884.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
334.0000000000,15827.,1225.6,3210.8,3490.4,2038.8,2355.6,6432.0,1114.5,2972.1,533.49,1180.1,1426.2,0.0000,-4421.3,-7297.0,-396.76,-3280.8,-3176.4,-14343.,-1733.3,-1525.9,-5396.9,-3083.1,-5882.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
335.0000000000,15838.,1219.2,3210.9,3414.3,2023.7,2334.1,6426.1,1114.6,2929.3,532.54,1186.3,1417.6,0.0000,-4411.9,-7286.8,-395.61,-3278.8,-3172.7,-14341.,-1732.4,-1521.9,-5395.7,-3082.7,-5880.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
336.0000000000,15834.,1226.0,3215.9,3412.2,2015.7,2286.2,6423.2,1112.9,2895.1,533.70,1177.4,1413.8,0.0000,-4402.9,-7278.6,-394.61,-3276.9,-3169.1,-14338.,-1731.8,-1518.3,-5395.0,-3082.1,-5878.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
337.0000000000,15824.,1232.0,3223.1,3405.2,2017.0,2280.1,6379.7,1119.7,2853.3,535.79,1164.9,1410.0,0.0000,-4394.4,-7270.7,-393.73,-3275.3,-3165.7,-14334.,-1731.3,-1515.0,-5394.1,-3081.6,-5877.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
338.0000000000,15314.,1233.3,3217.0,3378.0,1985.7,2276.2,6356.8,1122.4,2830.4,536.86,1135.6,1400.0,0.0000,-4386.5,-7263.3,-392.92,-3273.5,-3162.2,-14331.,-1730.9,-1512.0,-5393.5,-3081.5,-5876.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
339.0000000000,15198.,1229.1,3211.7,3375.4,1977.8,2277.7,6213.5,1118.7,2741.3,534.40,1116.1,1394.8,0.0000,-4378.7,-7256.2,-392.17,-3271.6,-3158.9,-14328.,-1730.6,-1509.2,-5393.0,-3081.1,-5874.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
340.0000000000,15193.,1230.4,3010.5,3379.4,1973.6,2298.6,6209.1,1108.4,2729.6,532.00,1104.6,1389.6,0.0000,-4420.4,-7274.7,-395.68,-3270.1,-3184.0,-14325.,-1732.0,-1534.9,-5404.3,-3083.3,-5882.3,11156.,4986.3,3819.7,3584.9,6949.4,2394.7,8583.9,2480.5,3792.1,1131.9,1626.7,1959.5,0.0000,-13.100,-13.884,-1.8060,-11.666,-10.733,-45.058,-35.642,-3.6120,-32.091,-4.3278,-44.141
341.0000000000,15192.,1209.3,2609.9,3371.4,1973.7,2295.9,6210.9,1102.3,2715.0,531.00,1094.0,1383.8,0.0000,-4389.9,-7270.0,-394.73,-3268.4,-3163.5,-14322.,-1731.4,-1519.8,-5395.9,-3081.6,-5876.2,40.576,18.137,13.893,13.039,25.277,8.7104,31.222,9.0224,13.793,4.1171,5.9169,7.1273,0.0000,-0.47601E-01,-0.50476E-01,-0.65689E-02,-0.42400E-01,-0.38968E-01,-0.16385,-0.12963,-0.13138E-01,-0.11672,-0.15739E-01,-0.16055
342.0000000000,15118.,1215.4,2615.9,3370.9,1948.7,2289.3,6186.8,1101.2,2707.4,530.37,1080.5,1375.7,0.0000,-4378.3,-7261.0,-393.34,-3266.5,-3158.3,-14319.,-1730.9,-1513.7,-5393.3,-3080.9,-5873.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
343.0000000000,15048.,1207.1,2621.1,3370.7,1950.4,2288.6,6108.9,1099.6,2707.5,529.44,1068.3,1366.5,0.0000,-4369.3,-7251.9,-392.11,-3264.6,-3154.5,-14315.,-1730.5,-1509.6,-5392.0,-3080.4,-5872.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
344.0000000000,15052.,1202.9,2621.6,3334.4,1933.6,2289.3,6087.9,1093.0,2686.3,527.61,1058.1,1359.8,0.0000,-4361.0,-7243.4,-391.08,-3262.6,-3151.1,-14313.,-1730.2,-1506.1,-5391.0,-3080.1,-5870.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
345.0000000000,15002.,1201.1,2597.4,3334.9,1927.2,2280.0,6081.7,1089.8,2677.2,527.02,1055.8,1349.0,0.0000,-4353.2,-7235.8,-390.19,-3260.6,-3147.9,-14310.,-1729.9,-1503.0,-5390.0,-3079.6,-5869.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
346.0000000000,14839.,1202.2,2574.0,3319.2,1895.1,2276.9,6047.6,1086.4,2671.6,527.44,1055.0,1349.1,0.0000,-4346.0,-7228.9,-389.41,-3258.7,-3145.0,-14306.,-1729.7,-1500.2,-5389.2,-3079.2,-5867.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
347.0000000000,14811.,1181.3,2564.9,3267.4,1899.8,2266.4,6016.4,1080.0,2669.0,527.69,1039.2,1349.7,0.0000,-4339.0,-7222.3,-388.69,-3256.7,-3142.0,-14303.,-1729.5,-1497.5,-5388.5,-3078.8,-5866.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
348.0000000000,14795.,1168.8,2557.5,3256.8,1907.2,2259.2,6014.2,1074.3,2667.6,524.98,1033.2,1348.9,0.0000,-4332.2,-7216.2,-388.02,-3254.8,-3139.1,-14299.,-1729.4,-1495.0,-5387.8,-3078.4,-5865.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
349.0000000000,14778.,1177.7,2559.0,3153.0,1924.2,2242.9,5991.9,1066.7,2667.7,518.02,1028.4,1337.0,0.0000,-4325.8,-7210.4,-387.38,-3252.9,-3136.2,-14296.,-1729.2,-1492.4,-5387.2,-3077.8,-5864.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
350.0000000000,14635.,1172.7,2557.7,3128.8,1915.0,2245.6,5979.8,1067.6,2676.7,521.00,1010.1,1320.3,0.0000,-4319.5,-7204.8,-386.76,-3251.0,-3133.4,-14293.,-1729.0,-1489.9,-5386.5,-3077.1,-5864.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
351.0000000000,14625.,1155.5,2553.3,3087.9,1884.4,2252.5,5951.8,1069.2,2686.4,522.06,1006.8,1312.6,0.0000,-4313.2,-7199.5,-386.16,-3249.2,-3130.6,-14291.,-1728.9,-1487.6,-5385.8,-3076.4,-5863.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
352.0000000000,14622.,1158.5,2553.4,3054.2,1853.4,2254.8,5968.8,1069.1,2629.7,521.92,1004.4,1310.8,0.0000,-4307.2,-7194.4,-385.58,-3247.3,-3127.8,-14289.,-1728.8,-1485.5,-5385.1,-3075.7,-5862.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
353.0000000000,14572.,1153.1,2556.9,3002.2,1847.4,2265.8,5947.5,1068.2,2609.5,519.76,1000.8,1298.9,0.0000,-4301.4,-7189.7,-385.00,-3245.5,-3125.1,-14288.,-1728.6,-1483.5,-5384.6,-3074.9,-5861.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
354.0000000000,14270.,1166.0,2554.3,2990.1,1845.4,2261.8,5927.6,1068.7,2605.2,518.81,999.02,1296.2,0.0000,-4295.8,-7185.0,-384.45,-3243.7,-3122.5,-14286.,-1728.5,-1481.7,-5384.1,-3074.2,-5860.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
355.0000000000,13915.,1172.1,2556.0,2978.7,1834.1,2266.5,5863.6,1069.4,2595.5,518.93,979.12,1287.7,0.0000,-4339.0,-7204.8,-388.10,-3242.3,-3148.1,-14284.,-1734.3,-1507.6,-5396.3,-3076.2,-5868.8,43056.,19245.,14742.,13836.,26822.,9242.7,33130.,9573.8,14636.,4368.7,6278.5,7562.8,0.0000,-49.942,-53.100,-6.9704,-44.720,-40.639,-173.39,-137.44,-13.941,-123.73,-16.651,-170.31
356.0000000000,13886.,1185.6,2554.8,2942.0,1818.3,2274.0,5849.8,1068.3,2579.7,517.70,972.84,1289.0,0.0000,-4359.5,-7227.0,-391.48,-3241.1,-3156.5,-14281.,-1735.0,-1522.2,-5400.4,-3076.8,-5871.9,16211.,7246.2,5550.8,5209.6,10099.,3480.1,12474.,3604.7,5510.8,1644.9,2364.0,2847.6,0.0000,-18.838,-20.010,-2.6245,-16.853,-15.321,-65.275,-51.748,-5.2490,-46.585,-6.2690,-64.126
357.0000000000,13859.,1167.6,2549.5,2935.9,1817.9,2219.5,5805.5,1068.5,2572.6,514.80,973.32,1292.4,0.0000,-4326.6,-7222.7,-389.89,-3239.6,-3134.3,-14277.,-1733.2,-1504.6,-5390.1,-3074.3,-5864.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
358.0000000000,13475.,1141.3,2542.9,2938.3,1789.6,2222.6,5756.3,1066.9,2521.7,509.74,974.75,1285.3,0.0000,-4314.6,-7214.3,-387.99,-3238.0,-3128.6,-14274.,-1731.7,-1497.5,-5386.6,-3073.2,-5861.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
359.0000000000,13126.,1134.0,2535.1,2933.1,1789.4,2217.7,5680.9,1067.6,2484.8,509.67,963.34,1261.1,0.0000,-4305.4,-7205.7,-386.40,-3236.3,-3124.8,-14272.,-1730.6,-1492.9,-5384.8,-3072.3,-5859.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
360.0000000000,13122.,1104.1,2550.7,2939.5,1829.9,2230.2,5662.5,1066.1,2488.7,505.20,959.93,1260.1,0.0000,-4346.3,-7222.2,-389.32,-3234.6,-3149.7,-14270.,-1731.7,-1517.1,-5395.5,-3074.4,-5866.2,14278.,6382.0,4888.8,4588.3,8894.6,3065.0,10986.,3174.8,4853.5,1448.7,2082.1,2508.0,0.0000,-16.570,-17.603,-2.3115,-14.826,-13.443,-57.460,-45.567,-4.6230,-41.018,-5.5174,-56.476
361.0000000000,13105.,1089.6,2558.4,2927.1,1829.1,2223.7,5654.2,1065.7,2498.9,505.85,960.00,1250.2,0.0000,-4365.0,-7241.3,-392.19,-3233.0,-3157.7,-14268.,-1734.6,-1529.9,-5399.1,-3075.2,-5868.9,28875.,12907.,9886.8,9279.1,17988.,6198.6,22219.,6420.6,9815.6,2929.8,4210.7,5072.0,0.0000,-33.565,-35.627,-4.6746,-30.008,-27.217,-116.19,-92.150,-9.3493,-82.949,-11.157,-114.21
362.0000000000,13070.,1081.6,2557.0,2924.3,1790.1,2188.2,5573.9,1063.8,2499.1,504.97,957.50,1238.8,0.0000,-4379.7,-7259.4,-394.46,-3231.5,-3163.6,-14265.,-1736.2,-1539.2,-5400.9,-3075.6,-5870.4,25096.,11218.,8592.9,8064.8,15634.,5387.4,19311.,5580.3,8531.0,2546.4,3659.6,4408.2,0.0000,-29.220,-30.990,-4.0629,-26.099,-23.677,-100.97,-80.089,-8.1257,-72.090,-9.6963,-99.269
363.0000000000,12809.,1077.0,2548.7,2917.3,1785.3,2166.3,5551.2,1064.4,2499.3,505.72,947.29,1228.4,0.0000,-4343.3,-7250.8,-392.01,-3229.7,-3140.4,-14261.,-1733.9,-1518.2,-5389.6,-3073.1,-5862.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
364.0000000000,12683.,1082.0,2551.8,2900.4,1797.4,2155.6,5537.2,1070.5,2464.9,506.76,936.42,1224.8,0.0000,-4328.9,-7238.5,-389.48,-3227.8,-3134.1,-14256.,-1732.1,-1509.1,-5385.8,-3071.9,-5859.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
365.0000000000,12008.,1068.2,2550.7,2901.7,1799.0,2151.1,5537.6,1060.4,2446.1,500.49,932.31,1223.9,0.0000,-4318.0,-7226.3,-387.45,-3225.8,-3129.9,-14252.,-1730.7,-1503.0,-5383.7,-3071.0,-5856.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
366.0000000000,11929.,1062.2,2560.6,2899.3,1815.7,2153.2,5508.3,1060.3,2448.0,497.41,934.52,1212.7,0.0000,-4308.6,-7215.2,-385.86,-3224.2,-3126.3,-14249.,-1729.7,-1498.1,-5382.4,-3070.3,-5854.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
367.0000000000,11855.,1070.1,2559.3,2897.2,1812.1,2153.4,5508.3,1060.5,2448.3,497.90,937.85,1206.9,0.0000,-4300.6,-7205.2,-384.59,-3222.4,-3123.1,-14246.,-1728.9,-1493.9,-5381.2,-3069.9,-5853.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
368.0000000000,11617.,1065.9,2558.8,2889.3,1805.5,2137.8,5473.6,1058.3,2449.1,498.96,932.94,1203.1,0.0000,-4293.2,-7196.9,-383.54,-3220.4,-3119.9,-14243.,-1728.3,-1490.1,-5380.3,-3069.5,-5851.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
369.0000000000,11001.,1074.3,2554.8,2841.7,1797.9,2134.9,5436.7,1046.1,2425.8,498.62,930.68,1200.7,0.0000,-4286.0,-7189.2,-382.64,-3218.7,-3116.7,-14240.,-1727.9,-1486.7,-5379.7,-3069.2,-5850.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
370.0000000000,10961.,1074.9,2553.0,2815.8,1770.8,2128.1,5333.5,1045.4,2411.5,498.70,921.02,1203.7,0.0000,-4279.0,-7182.0,-381.84,-3216.9,-3113.5,-14237.,-1727.5,-1483.5,-5379.5,-3068.8,-5849.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
371.0000000000,10903.,1076.1,2553.3,2806.3,1771.0,2128.9,5304.1,1042.1,2407.7,492.72,914.26,1195.7,0.0000,-4272.1,-7175.3,-381.11,-3215.0,-3110.3,-14234.,-1727.3,-1480.7,-5378.9,-3068.0,-5848.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
372.0000000000,10902.,1078.8,2554.0,2806.4,1738.8,2119.7,5270.5,1042.6,2408.4,488.06,908.04,1194.2,0.0000,-4265.4,-7168.9,-380.42,-3213.3,-3107.3,-14231.,-1727.0,-1478.1,-5378.3,-3067.3,-5847.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
373.0000000000,10382.,1063.7,2540.3,2782.2,1688.2,2117.9,5220.9,1034.2,2426.8,486.88,907.11,1196.5,0.0000,-4259.5,-7161.9,-379.78,-3211.8,-3104.4,-14229.,-1726.8,-1475.7,-5377.6,-3066.7,-5846.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
374.0000000000,10125.,1065.5,2531.2,2771.4,1672.1,2118.1,5103.5,1022.8,2429.6,487.08,910.08,1194.6,0.0000,-4253.7,-7155.4,-379.17,-3210.2,-3101.6,-14226.,-1726.6,-1473.4,-5377.0,-3066.3,-5845.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
375.0000000000,10121.,1081.5,2533.4,2772.4,1648.6,2118.4,5057.0,1021.7,2435.6,486.56,905.28,1183.0,0.0000,-4248.0,-7149.5,-378.59,-3208.5,-3098.8,-14223.,-1726.5,-1471.3,-5376.5,-3065.9,-5844.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
376.0000000000,10103.,1091.6,2528.0,2769.7,1650.1,2109.1,4919.0,1016.7,2401.8,485.69,896.27,1170.3,0.0000,-4242.2,-7144.2,-378.01,-3206.7,-3095.8,-14220.,-1726.3,-1469.2,-5376.0,-3065.2,-5844.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
377.0000000000,10075.,1093.9,2520.5,2771.5,1658.1,2114.7,4833.1,1016.9,2371.7,485.00,898.29,1170.1,0.0000,-4236.6,-7139.3,-377.46,-3205.2,-3093.1,-14217.,-1726.1,-1467.3,-5375.4,-3064.6,-5843.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
378.0000000000,10092.,1095.3,2514.7,2730.8,1654.2,2123.0,4806.5,1013.2,2352.3,484.16,899.18,1168.1,0.0000,-4230.8,-7134.5,-376.92,-3203.6,-3090.2,-14215.,-1726.0,-1465.4,-5374.9,-3064.0,-5842.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
379.0000000000,10105.,1102.1,2517.5,2728.2,1658.1,2123.8,4768.0,1005.5,2343.9,485.23,899.99,1168.7,0.0000,-4225.2,-7129.9,-376.39,-3201.9,-3087.4,-14212.,-1725.9,-1463.7,-5374.5,-3063.7,-5842.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
380.0000000000,10078.,1109.0,2512.7,2723.9,1658.8,2122.2,4688.3,986.92,2339.2,483.42,889.68,1170.7,0.0000,-4219.8,-7125.7,-375.89,-3200.2,-3084.7,-14209.,-1725.7,-1462.0,-5374.0,-3063.4,-5841.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
381.0000000000,10063.,1102.8,2519.4,2716.7,1635.4,2123.1,4623.9,983.59,2342.5,481.32,881.63,1170.1,0.0000,-4214.6,-7121.6,-375.38,-3198.5,-3082.1,-14207.,-1725.6,-1460.3,-5373.4,-3063.0,-5840.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
382.0000000000,10048.,1095.5,2525.0,2645.5,1620.2,2084.0,4571.5,974.77,2342.2,480.71,876.06,1150.2,0.0000,-4209.4,-7117.6,-374.89,-3196.8,-3079.5,-14204.,-1725.5,-1458.7,-5372.9,-3062.6,-5840.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
383.0000000000,9851.6,1098.1,2526.9,2614.2,1622.9,2064.5,4559.4,974.64,2344.0,479.54,876.68,1147.2,0.0000,-4204.3,-7113.8,-374.41,-3195.1,-3077.0,-14202.,-1725.3,-1457.1,-5372.5,-3062.2,-5839.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
384.0000000000,9789.3,1120.8,2526.5,2613.7,1618.7,2032.3,4534.5,975.25,2344.1,480.82,871.48,1142.7,0.0000,-4199.3,-7110.1,-373.93,-3193.4,-3074.5,-14199.,-1725.2,-1455.5,-5372.1,-3061.8,-5838.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
385.0000000000,9744.8,1123.6,2529.3,2617.2,1596.1,2011.0,4527.2,973.08,2301.3,481.46,856.93,1139.2,0.0000,-4194.3,-7106.3,-373.45,-3191.8,-3072.1,-14197.,-1725.1,-1454.0,-5371.7,-3061.5,-5838.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
386.0000000000,9731.1,1123.6,2533.2,2607.5,1602.0,2007.4,4508.2,967.97,2298.7,480.79,847.89,1138.8,0.0000,-4189.4,-7102.6,-372.98,-3190.1,-3069.7,-14194.,-1725.0,-1452.5,-5371.4,-3061.2,-5837.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
387.0000000000,9727.0,1126.8,2533.8,2540.5,1599.6,2011.4,4488.0,959.94,2298.2,481.08,846.44,1121.4,0.0000,-4184.5,-7099.4,-372.52,-3188.4,-3067.3,-14192.,-1724.9,-1451.1,-5371.1,-3060.8,-5836.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
388.0000000000,9727.1,1127.9,2530.5,2509.3,1600.4,2015.1,4463.4,960.30,2294.9,482.20,834.66,1120.3,0.0000,-4179.8,-7096.5,-372.06,-3186.6,-3064.9,-14189.,-1724.7,-1449.8,-5370.8,-3060.3,-5836.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
389.0000000000,9716.4,1139.9,2538.8,2449.3,1597.4,2006.8,4450.0,959.49,2297.6,482.89,830.06,1104.9,0.0000,-4223.2,-7117.3,-375.78,-3185.2,-3090.8,-14188.,-1725.2,-1475.1,-5382.1,-3062.6,-5843.9,3723.5,1664.3,1274.9,1196.6,2319.6,799.32,2865.1,827.95,1265.7,377.81,542.98,654.04,0.0000,-4.2425,-4.5197,-0.60280,-3.8291,-3.3878,-14.943,-11.869,-1.2056,-10.683,-1.4304,-14.740
390.0000000000,9682.3,1142.7,2538.6,2434.1,1596.7,1981.8,4459.9,959.90,2287.0,484.05,822.84,1086.1,0.0000,-4195.9,-7116.1,-375.05,-3183.7,-3071.3,-14185.,-1725.0,-1462.4,-5373.9,-3060.6,-5838.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
391.0000000000,9645.0,1139.0,2524.6,2431.5,1603.4,1968.0,4460.8,960.57,2285.8,484.21,817.43,1081.8,0.0000,-4187.2,-7111.1,-373.85,-3182.1,-3066.7,-14182.,-1724.7,-1457.6,-5371.5,-3059.8,-5836.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
392.0000000000,9489.2,1134.0,2526.2,2410.7,1605.9,1968.7,4461.7,959.08,2258.9,474.40,816.38,1076.6,0.0000,-4180.7,-7105.8,-372.78,-3180.5,-3063.6,-14179.,-1724.5,-1454.6,-5370.4,-3059.1,-5834.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
393.0000000000,9498.9,1132.2,2424.8,2389.6,1603.8,1978.0,4465.8,956.32,2231.8,467.18,806.31,1063.2,0.0000,-4174.9,-7100.7,-371.89,-3178.9,-3060.9,-14177.,-1724.3,-1452.3,-5369.6,-3058.5,-5834.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
394.0000000000,9389.4,1128.8,1911.6,2353.7,1606.6,1980.6,4480.9,957.68,2210.6,463.35,803.69,1063.1,0.0000,-4169.6,-7095.9,-371.14,-3177.3,-3058.4,-14174.,-1724.2,-1450.2,-5369.1,-3057.9,-5833.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
395.0000000000,9374.6,1126.1,1912.6,2353.4,1607.6,1977.9,4481.3,958.33,2184.9,463.51,798.16,1055.9,0.0000,-4164.5,-7091.3,-370.48,-3175.7,-3056.0,-14171.,-1724.0,-1448.3,-5368.5,-3057.3,-5832.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
396.0000000000,9334.9,1123.2,1912.7,2326.2,1611.6,1976.1,4463.5,958.59,2181.3,456.65,793.82,1039.4,0.0000,-4159.6,-7087.0,-369.88,-3174.2,-3053.6,-14168.,-1723.9,-1446.6,-5368.1,-3056.7,-5831.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
397.0000000000,9259.1,1134.2,1912.1,2314.4,1613.6,1969.7,4427.9,958.41,2183.3,453.14,785.82,1034.7,0.0000,-4155.0,-7083.1,-369.32,-3172.7,-3051.3,-14166.,-1723.7,-1444.9,-5367.6,-3056.2,-5830.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
398.0000000000,9168.8,1139.8,1913.1,2325.0,1614.9,1968.1,4378.4,954.56,2178.8,453.68,784.66,1033.2,0.0000,-4150.3,-7079.4,-368.81,-3171.1,-3049.0,-14163.,-1723.6,-1443.2,-5367.2,-3055.7,-5830.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
399.0000000000,9145.6,1142.9,1911.4,2318.9,1610.2,1958.9,4341.4,941.03,2167.9,452.11,778.02,1025.9,0.0000,-4145.6,-7075.8,-368.29,-3169.6,-3046.6,-14160.,-1723.5,-1441.5,-5366.9,-3055.2,-5829.3,127.82,57.134,43.766,41.076,79.628,27.439,98.355,28.422,43.451,12.969,18.639,22.452,0.0000,-0.14452,-0.15411,-0.20693E-01,-0.13087,-0.11466,-0.51239,-0.40723,-0.41386E-01,-0.36659,-0.48989E-01,-0.50602
400.0000000000,9145.7,1143.6,1912.3,2318.5,1605.7,1948.2,4335.2,927.23,2157.1,446.56,776.34,1021.2,0.0000,-4141.1,-7072.5,-367.77,-3168.0,-3044.2,-14158.,-1723.4,-1440.0,-5366.6,-3054.6,-5828.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
401.0000000000,9158.4,1148.4,1913.5,2321.4,1612.8,1948.6,4318.7,924.21,2144.0,447.35,777.73,1016.7,0.0000,-4136.8,-7069.4,-367.27,-3166.5,-3042.0,-14155.,-1723.2,-1438.5,-5366.3,-3054.1,-5828.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
402.0000000000,9117.6,1141.8,1917.4,2317.5,1611.2,1958.3,4302.0,917.67,2140.6,446.77,768.85,1018.6,0.0000,-4132.7,-7066.2,-366.78,-3164.9,-3039.7,-14152.,-1723.1,-1437.1,-5366.0,-3053.6,-5827.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
403.0000000000,8763.4,1137.3,1927.4,2317.9,1615.4,1956.1,4299.7,918.91,2142.4,445.97,766.86,1007.9,0.0000,-4128.7,-7063.2,-366.30,-3163.4,-3037.4,-14149.,-1723.0,-1435.7,-5365.7,-3053.1,-5826.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
404.0000000000,8534.8,1127.8,1930.8,2285.4,1618.6,1948.0,4297.4,916.73,2140.6,448.35,760.90,1009.7,0.0000,-4124.7,-7060.2,-365.84,-3161.9,-3035.2,-14146.,-1722.9,-1434.3,-5365.4,-3052.6,-5826.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
405.0000000000,8544.1,1127.2,1931.1,2275.5,1614.9,1944.7,4261.1,909.03,2147.6,448.61,755.27,1009.9,0.0000,-4120.7,-7057.0,-365.38,-3160.3,-3033.0,-14143.,-1722.8,-1433.1,-5365.2,-3052.2,-5825.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
406.0000000000,8549.1,1126.5,1932.5,2274.1,1620.5,1913.3,4184.5,906.14,2127.6,448.12,756.46,1005.7,0.0000,-4116.8,-7053.9,-364.95,-3158.8,-3030.8,-14141.,-1722.7,-1431.8,-5365.0,-3051.7,-5824.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
407.0000000000,8416.3,1117.6,1933.2,2269.7,1617.7,1901.5,4129.5,903.09,2106.6,444.82,756.64,1000.9,0.0000,-4112.8,-7050.9,-364.51,-3157.2,-3028.5,-14138.,-1722.5,-1430.7,-5364.7,-3051.3,-5823.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
408.0000000000,8321.5,1108.8,1933.9,2266.0,1618.0,1901.3,4097.3,894.73,2074.0,440.56,755.56,1001.6,0.0000,-4108.9,-7048.0,-364.08,-3155.6,-3026.4,-14136.,-1722.4,-1429.5,-5364.5,-3050.8,-5823.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
409.0000000000,8317.3,1111.7,1935.2,2218.6,1583.8,1902.2,4100.1,896.45,2072.9,437.89,750.42,998.35,0.0000,-4105.0,-7045.4,-363.66,-3154.0,-3024.2,-14133.,-1722.3,-1428.4,-5364.1,-3050.4,-5822.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
410.0000000000,8306.8,1111.4,1938.4,2144.6,1583.5,1890.6,4110.1,896.05,2049.7,437.46,752.22,987.07,0.0000,-4101.1,-7042.8,-363.25,-3152.5,-3022.1,-14131.,-1722.2,-1427.3,-5363.8,-3049.9,-5821.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
411.0000000000,8307.3,1108.3,1936.2,2140.5,1572.8,1872.2,4106.6,897.90,2035.0,436.72,753.74,983.37,0.0000,-4097.4,-7040.3,-362.84,-3150.9,-3020.0,-14129.,-1722.1,-1426.3,-5363.5,-3049.4,-5820.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
412.0000000000,8317.4,1108.6,1935.4,2113.9,1547.6,1870.0,4098.4,896.49,2031.8,435.36,755.47,984.72,0.0000,-4093.6,-7037.8,-362.43,-3149.4,-3018.0,-14126.,-1722.0,-1425.3,-5363.1,-3049.0,-5820.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
413.0000000000,8240.1,1111.1,1935.5,2101.6,1535.2,1869.6,4004.3,878.40,2032.7,434.22,747.28,973.68,0.0000,-4089.9,-7035.4,-362.03,-3147.9,-3015.9,-14124.,-1721.8,-1424.3,-5362.7,-3048.5,-5819.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
414.0000000000,8136.6,1107.8,1931.8,2101.9,1525.6,1833.2,3984.2,870.27,2030.3,434.86,740.57,971.68,0.0000,-4086.2,-7033.0,-361.63,-3146.4,-3013.8,-14122.,-1721.7,-1423.4,-5362.4,-3048.0,-5819.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
415.0000000000,8090.2,1108.9,1924.5,2072.9,1525.8,1832.3,3983.4,871.26,2033.3,435.75,742.18,972.89,0.0000,-4082.5,-7030.6,-361.23,-3144.9,-3011.8,-14120.,-1721.6,-1422.4,-5362.0,-3047.5,-5818.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
416.0000000000,7940.9,1112.2,1920.8,2071.3,1532.1,1825.8,3983.6,874.25,2036.7,437.22,743.16,974.93,0.0000,-4078.9,-7028.4,-360.83,-3143.3,-3009.8,-14118.,-1721.5,-1421.5,-5361.6,-3047.1,-5818.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
417.0000000000,7938.5,1116.9,1919.8,2071.9,1540.1,1823.3,3958.0,873.34,2037.5,438.55,726.78,969.68,0.0000,-4075.3,-7026.1,-360.45,-3141.8,-3007.8,-14116.,-1721.4,-1420.6,-5361.3,-3046.6,-5817.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
418.0000000000,7963.8,1119.2,1919.5,2072.2,1542.0,1808.7,3958.3,865.85,2033.1,438.54,724.31,959.97,0.0000,-4071.7,-7024.0,-360.07,-3140.3,-3005.8,-14114.,-1721.3,-1419.7,-5360.9,-3046.2,-5816.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
419.0000000000,7945.8,1122.2,1945.0,2072.1,1549.3,1788.2,3960.2,866.12,2021.9,439.10,718.08,960.96,0.0000,-4068.1,-7021.9,-359.70,-3138.8,-3003.8,-14112.,-1721.1,-1418.9,-5360.5,-3045.8,-5816.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
420.0000000000,7884.2,1115.6,1942.8,2059.1,1547.4,1785.6,3928.6,860.03,2020.0,439.86,713.25,955.58,0.0000,-4064.6,-7019.7,-359.33,-3137.4,-3001.8,-14109.,-1721.0,-1418.1,-5360.1,-3045.3,-5815.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
421.0000000000,7826.7,1105.3,1951.5,2022.6,1548.4,1797.3,3891.5,847.12,2025.0,439.18,706.24,954.92,0.0000,-4108.3,-7041.1,-363.12,-3136.2,-3028.0,-14108.,-1721.3,-1443.0,-5371.4,-3047.6,-5823.0,2550.5,1140.0,873.28,819.60,1588.8,547.50,1962.5,567.11,866.98,258.78,371.92,447.99,0.0000,-2.8499,-3.0304,-0.41290,-2.5951,-2.2318,-10.200,-8.1167,-0.82579,-7.3074,-0.97209,-10.096
422.0000000000,7808.0,1102.9,1954.9,2027.8,1539.5,1768.2,3883.5,850.47,2025.3,438.84,706.56,954.88,0.0000,-4129.8,-7064.3,-366.66,-3135.2,-3037.1,-14107.,-1726.3,-1457.8,-5375.7,-3048.3,-5826.6,37393.,16714.,12803.,12016.,23294.,8026.9,28772.,8314.5,12711.,3794.0,5452.7,6568.1,0.0000,-41.872,-44.478,-6.0535,-38.086,-32.771,-149.54,-119.00,-12.107,-107.13,-14.250,-148.02
423.0000000000,7792.8,1103.2,1956.8,2021.0,1537.8,1771.8,3875.1,852.24,2036.6,437.01,708.84,956.68,0.0000,-4147.2,-7085.5,-369.47,-3134.3,-3043.9,-14105.,-1726.5,-1469.1,-5377.8,-3048.7,-5828.3,11449.,5117.7,3920.3,3679.3,7132.5,2457.8,8809.9,2545.9,3892.0,1161.7,1669.6,2011.1,0.0000,-12.848,-13.636,-1.8536,-11.672,-10.047,-45.785,-36.436,-3.7071,-32.802,-4.3625,-45.324
424.0000000000,7727.3,1098.1,1953.3,2015.7,1538.0,1714.4,3832.0,848.39,2031.7,437.43,710.63,955.84,0.0000,-4114.7,-7080.5,-367.48,-3133.1,-3021.7,-14102.,-1724.9,-1451.4,-5366.9,-3046.2,-5820.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
425.0000000000,7592.4,1094.2,1953.4,2002.0,1553.8,1684.9,3826.0,844.86,2020.6,430.21,712.31,953.93,0.0000,-4103.6,-7071.8,-365.33,-3131.6,-3016.1,-14100.,-1723.7,-1444.1,-5363.4,-3045.0,-5817.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
426.0000000000,7438.9,1074.9,1944.5,1987.5,1622.8,1673.2,3829.7,831.46,2020.5,427.89,712.27,950.58,0.0000,-4095.7,-7063.2,-363.61,-3130.1,-3012.5,-14098.,-1722.8,-1439.5,-5361.6,-3044.2,-5815.9,1054.2,471.21,360.96,338.77,656.73,226.30,811.18,234.41,358.36,106.97,153.73,185.17,0.0000,-1.1801,-1.2541,-0.17067,-1.0725,-0.91995,-4.2149,-3.3545,-0.34133,-3.0198,-0.40132,-4.1733
427.0000000000,7439.6,1066.8,1956.7,1988.1,1679.2,1656.9,3829.5,824.49,2014.7,428.22,711.27,940.82,0.0000,-4089.0,-7055.6,-362.28,-3128.5,-3009.4,-14096.,-1722.1,-1435.9,-5360.5,-3043.5,-5814.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
428.0000000000,7339.0,1064.2,1958.3,1989.1,1677.8,1652.6,3817.2,817.01,1990.4,428.04,709.24,940.23,0.0000,-4083.0,-7048.9,-361.25,-3126.9,-3006.6,-14094.,-1721.5,-1432.8,-5359.5,-3042.8,-5813.3,107.44,48.025,36.788,34.527,66.932,23.064,82.673,23.891,36.523,10.902,15.668,18.872,0.0000,-0.12007,-0.12761,-0.17394E-01,-0.10920,-0.93477E-01,-0.42952,-0.34185,-0.34788E-01,-0.30774,-0.40878E-01,-0.42533
429.0000000000,7263.7,1068.2,1940.1,1989.9,1668.5,1651.4,3783.1,815.74,1988.6,426.96,693.55,939.87,0.0000,-4077.5,-7043.0,-360.41,-3125.4,-3004.0,-14092.,-1721.0,-1429.9,-5358.8,-3042.0,-5812.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
430.0000000000,7235.9,1062.5,1938.6,1975.9,1669.6,1649.7,3756.1,806.94,1961.1,425.90,687.67,938.19,0.0000,-4072.3,-7037.6,-359.71,-3124.0,-3001.4,-14090.,-1720.7,-1427.3,-5357.9,-3041.3,-5811.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
431.0000000000,7237.9,1058.0,1943.3,1948.1,1676.8,1656.2,3715.8,806.13,1959.4,426.73,688.81,933.43,0.0000,-4067.4,-7032.7,-359.11,-3122.5,-2998.8,-14088.,-1720.4,-1425.2,-5357.2,-3040.7,-5810.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
432.0000000000,7234.3,1060.2,1942.8,1942.4,1678.1,1659.9,3671.1,806.63,1962.8,427.06,685.43,924.85,0.0000,-4062.8,-7028.0,-358.57,-3121.1,-2996.3,-14087.,-1720.2,-1423.3,-5356.5,-3040.1,-5809.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
433.0000000000,7229.6,1056.7,1945.0,1946.8,1680.4,1661.4,3652.8,807.22,1926.4,426.97,681.54,915.68,0.0000,-4058.3,-7023.9,-358.09,-3119.7,-2993.9,-14085.,-1720.0,-1421.5,-5355.8,-3039.5,-5808.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
434.0000000000,7212.2,1055.2,1956.2,1950.2,1683.9,1671.7,3650.0,803.21,1920.1,427.03,673.29,908.97,0.0000,-4101.2,-7043.4,-361.79,-3118.6,-3019.7,-14084.,-1720.1,-1445.9,-5366.7,-3041.6,-5816.3,1573.9,703.50,538.90,505.77,980.46,337.86,1211.1,349.97,535.01,159.69,229.51,276.46,0.0000,-1.7556,-1.8628,-0.25480,-1.5984,-1.3626,-6.2897,-5.0063,-0.50960,-4.5068,-0.59778,-6.2307
435.0000000000,7111.4,1051.2,1948.0,1944.5,1699.1,1661.5,3656.5,797.16,1919.2,423.90,673.60,906.57,0.0000,-4074.4,-7041.2,-361.10,-3117.4,-3000.1,-14082.,-1719.9,-1433.4,-5358.3,-3039.6,-5810.5,3.4756,1.5535,1.1901,1.1169,2.1652,0.74611,2.6744,0.77283,1.1815,0.35266,0.50683,0.61050,0.0000,-0.38746E-02,-0.41124E-02,-0.56267E-03,-0.35279E-02,-0.30038E-02,-0.13889E-01,-0.11055E-01,-0.11253E-02,-0.99519E-02,-0.13196E-02,-0.13759E-01
436.0000000000,7084.8,1055.6,1936.8,1929.8,1714.8,1648.3,3644.4,796.97,1914.3,423.48,675.07,894.33,0.0000,-4065.9,-7035.6,-359.95,-3116.1,-2995.4,-14081.,-1719.7,-1428.5,-5355.7,-3038.7,-5808.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
437.0000000000,7086.7,1068.0,1932.2,1900.9,1722.9,1608.4,3615.9,793.28,1902.6,424.73,667.73,888.74,0.0000,-4059.9,-7029.8,-358.95,-3114.8,-2992.3,-14079.,-1719.5,-1425.4,-5354.6,-3038.0,-5807.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
438.0000000000,6740.0,1070.1,1937.8,1900.1,1728.6,1619.7,3617.1,779.30,1895.6,425.41,667.39,876.29,0.0000,-4054.5,-7024.5,-358.13,-3113.4,-2989.5,-14077.,-1719.3,-1422.9,-5353.8,-3037.3,-5806.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
439.0000000000,6421.0,1068.9,1943.6,1897.0,1732.8,1626.0,3602.2,779.59,1900.9,425.08,669.00,875.12,0.0000,-4049.5,-7019.6,-357.45,-3112.1,-2986.8,-14076.,-1719.2,-1420.8,-5353.1,-3036.7,-5805.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
440.0000000000,6388.9,1062.7,1938.8,1892.2,1727.9,1627.6,3576.6,780.30,1900.8,423.09,667.23,876.05,0.0000,-4044.7,-7015.1,-356.87,-3110.7,-2984.3,-14074.,-1719.1,-1418.9,-5352.5,-3036.2,-5805.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
441.0000000000,6395.4,1064.6,1935.6,1852.5,1730.5,1629.0,3571.2,781.83,1898.8,423.91,662.19,877.83,0.0000,-4040.1,-7011.0,-356.36,-3109.3,-2981.8,-14073.,-1718.9,-1417.2,-5351.9,-3035.7,-5804.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
442.0000000000,6394.2,1074.0,1935.1,1853.0,1727.0,1609.8,3558.2,782.50,1889.8,423.91,662.69,869.65,0.0000,-4035.8,-7007.2,-355.90,-3107.8,-2979.3,-14071.,-1718.8,-1415.5,-5351.4,-3035.2,-5804.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
443.0000000000,6284.2,1075.5,1932.3,1858.1,1730.1,1577.1,3524.5,782.23,1875.9,423.12,663.53,869.93,0.0000,-4031.6,-7003.7,-355.47,-3106.2,-2976.9,-14070.,-1718.7,-1414.0,-5350.8,-3034.7,-5803.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
444.0000000000,6257.6,1080.1,1932.2,1829.6,1718.6,1525.9,3490.8,774.87,1855.0,422.97,666.41,864.19,0.0000,-4027.5,-7000.7,-355.07,-3104.6,-2974.5,-14069.,-1718.6,-1412.6,-5350.2,-3034.2,-5803.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
445.0000000000,6260.1,1096.9,1811.4,1777.8,1713.5,1472.2,3441.8,771.25,1835.9,420.29,667.53,862.37,0.0000,-4023.6,-6997.8,-354.69,-3103.1,-2972.2,-14067.,-1718.4,-1411.2,-5349.5,-3033.7,-5802.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
446.0000000000,6264.3,1097.1,1323.5,1744.9,1713.1,1450.4,3377.8,757.65,1829.8,413.25,669.93,863.08,0.0000,-4019.9,-6995.0,-354.32,-3101.6,-2969.8,-14066.,-1718.3,-1409.9,-5349.0,-3033.1,-5802.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
447.0000000000,6218.2,1096.8,1330.2,1727.0,1713.1,1442.1,3383.7,753.57,1836.0,413.45,671.83,864.47,0.0000,-4016.1,-6992.2,-353.96,-3100.1,-2967.4,-14065.,-1718.2,-1408.7,-5348.5,-3032.6,-5802.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
448.0000000000,6264.9,1100.9,1327.3,1715.6,1715.0,1455.5,3378.6,737.76,1842.3,412.52,671.57,856.80,0.0000,-4059.5,-7013.1,-357.75,-3099.0,-2993.3,-14064.,-1719.3,-1433.0,-5359.7,-3034.8,-5810.0,8387.8,3749.2,2872.0,2695.4,5225.2,1800.6,6454.1,1865.1,2851.3,851.06,1223.1,1473.3,0.0000,-9.2888,-9.8399,-1.3579,-8.4888,-7.1486,-33.504,-26.666,-2.7158,-24.004,-3.1730,-33.205
449.0000000000,6294.6,1089.4,1318.6,1719.9,1724.7,1436.4,3325.6,737.78,1839.0,411.07,671.50,855.55,0.0000,-4033.5,-7012.2,-357.15,-3097.7,-2973.8,-14062.,-1718.9,-1421.4,-5351.4,-3032.7,-5804.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
450.0000000000,6289.0,1086.0,1318.7,1719.7,1725.9,1402.7,3309.1,737.72,1849.0,410.01,669.32,848.35,0.0000,-4025.6,-7007.8,-356.07,-3096.3,-2969.3,-14060.,-1718.6,-1417.0,-5348.8,-3031.8,-5802.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
451.0000000000,6256.1,1090.4,1322.7,1728.0,1728.8,1414.2,3268.6,738.01,1864.8,410.55,662.00,846.81,0.0000,-4067.2,-7026.6,-359.27,-3095.3,-2994.4,-14059.,-1718.6,-1440.2,-5359.2,-3033.7,-5809.9,1438.8,643.12,492.65,462.37,896.32,308.87,1107.1,319.93,489.10,145.99,209.81,252.73,0.0000,-1.5945,-1.6875,-0.23293,-1.4564,-1.2244,-5.7465,-4.5738,-0.46586,-4.1171,-0.54389,-5.6957
452.0000000000,6261.4,1092.6,1315.6,1727.0,1722.9,1390.8,3231.9,737.89,1853.3,408.29,649.21,848.57,0.0000,-4039.8,-7023.4,-358.24,-3094.1,-2974.5,-14057.,-1718.3,-1427.3,-5350.5,-3031.5,-5804.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
453.0000000000,6216.9,1102.3,1314.6,1727.9,1720.4,1345.0,3192.0,737.47,1831.2,398.99,644.69,847.93,0.0000,-4031.0,-7017.1,-356.85,-3092.8,-2969.7,-14055.,-1718.0,-1422.1,-5347.8,-3030.5,-5802.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
454.0000000000,6235.4,1109.3,1311.8,1696.8,1721.4,1301.4,3200.5,739.98,1802.8,397.95,640.00,848.22,0.0000,-4024.7,-7010.7,-355.70,-3091.5,-2966.4,-14053.,-1717.8,-1418.8,-5346.4,-3029.7,-5801.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
455.0000000000,6239.9,1098.5,1319.0,1694.9,1721.6,1301.2,3184.7,726.47,1803.3,395.57,633.88,847.65,0.0000,-4019.2,-7004.8,-354.77,-3090.0,-2963.5,-14051.,-1717.6,-1416.2,-5345.4,-3029.0,-5800.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
456.0000000000,6194.4,1099.4,1323.3,1687.2,1721.7,1302.7,3153.1,721.92,1809.6,394.12,633.43,844.85,0.0000,-4014.2,-6999.3,-354.02,-3088.6,-2960.7,-14050.,-1717.5,-1413.9,-5344.7,-3028.3,-5800.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
457.0000000000,6165.5,1095.6,1323.8,1661.5,1724.0,1304.8,3136.5,712.94,1806.4,394.48,634.62,842.64,0.0000,-4009.4,-6994.2,-353.39,-3087.2,-2958.1,-14048.,-1717.3,-1411.9,-5344.0,-3027.6,-5799.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
458.0000000000,6132.4,1096.5,1328.0,1658.6,1724.3,1293.2,3119.7,713.18,1808.2,394.00,635.11,835.88,0.0000,-4004.9,-6989.6,-352.85,-3085.8,-2955.6,-14046.,-1717.2,-1410.1,-5343.4,-3026.9,-5799.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
459.0000000000,6079.8,1101.9,1343.2,1660.7,1725.0,1305.8,3113.6,695.26,1815.3,393.30,634.66,823.36,0.0000,-4047.5,-7008.9,-356.51,-3084.7,-2981.2,-14045.,-1721.4,-1433.9,-5355.1,-3028.9,-5807.7,31553.,14104.,10804.,10140.,19656.,6773.4,24279.,7016.1,10726.,3201.6,4601.2,5542.4,0.0000,-34.847,-36.851,-5.1082,-31.885,-26.628,-125.96,-100.28,-10.216,-90.256,-11.901,-124.88
460.0000000000,6032.3,1103.0,1355.6,1668.2,1727.3,1294.1,3070.2,679.36,1804.6,391.88,636.47,812.08,0.0000,-4020.9,-7006.8,-355.82,-3083.6,-2961.6,-14043.,-1720.2,-1421.8,-5347.0,-3026.8,-5802.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
461.0000000000,6027.7,1116.1,1364.5,1678.9,1732.2,1291.0,3016.8,677.55,1781.6,392.06,635.38,811.84,0.0000,-4059.7,-7024.9,-358.81,-3082.7,-2985.0,-14042.,-1719.5,-1442.8,-5355.9,-3028.4,-5808.9,1437.0,642.31,492.02,461.78,895.18,308.47,1105.7,319.53,488.48,145.80,209.55,252.41,0.0000,-1.5893,-1.6789,-0.23264,-1.4529,-1.2127,-5.7352,-4.5666,-0.46527,-4.1101,-0.54176,-5.6872
462.0000000000,5973.6,1114.1,1359.2,1671.5,1711.4,1273.6,2997.0,674.08,1748.8,392.20,634.78,814.26,0.0000,-4031.2,-7020.8,-357.55,-3081.6,-2964.6,-14040.,-1718.7,-1428.8,-5346.6,-3026.1,-5802.7,239.64,107.11,82.052,77.008,149.28,51.442,184.39,53.285,81.460,24.315,34.945,42.093,0.0000,-0.26486,-0.27991,-0.38795E-01,-0.24214,-0.20186,-0.95632,-0.76152,-0.77590E-01,-0.68539,-0.90319E-01,-0.94839
463.0000000000,5987.4,1120.9,1360.7,1648.0,1686.0,1249.3,3002.4,667.06,1722.9,391.45,638.31,805.62,0.0000,-4068.9,-7037.0,-360.15,-3080.7,-2987.6,-14039.,-1718.6,-1449.1,-5355.2,-3027.6,-5808.5,3497.5,1563.3,1197.5,1123.9,2178.8,750.79,2691.2,777.68,1188.9,354.87,510.01,614.33,0.0000,-3.8731,-4.0882,-0.56621,-3.5376,-2.9509,-13.956,-11.114,-1.1324,-10.003,-1.3180,-13.841
464.0000000000,6017.3,1117.8,1349.3,1632.3,1679.9,1240.4,3006.5,667.72,1704.8,382.97,639.49,805.03,0.0000,-4039.5,-7031.4,-358.60,-3079.6,-2966.9,-14037.,-1718.0,-1434.2,-5345.8,-3025.2,-5802.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
465.0000000000,5981.7,1116.0,1355.1,1637.6,1682.7,1220.7,3015.0,668.57,1684.7,376.19,638.28,793.04,0.0000,-4029.3,-7022.8,-356.84,-3078.4,-2961.5,-14035.,-1717.5,-1427.6,-5342.8,-3024.0,-5799.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
466.0000000000,5948.0,1113.0,1364.1,1636.6,1687.5,1204.0,2999.5,668.73,1690.0,373.35,628.13,784.65,0.0000,-4021.8,-7014.5,-355.41,-3077.1,-2957.9,-14033.,-1717.1,-1423.3,-5341.3,-3023.2,-5798.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
467.0000000000,5834.3,1113.7,1373.0,1638.6,1686.8,1204.8,2965.4,667.21,1689.1,368.57,622.11,776.60,0.0000,-4015.3,-7007.0,-354.29,-3075.7,-2954.7,-14032.,-1716.8,-1419.8,-5340.3,-3022.4,-5797.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
468.0000000000,5710.4,1113.0,1373.5,1639.4,1664.9,1203.8,2936.1,668.86,1655.8,358.53,613.49,776.28,0.0000,-4009.4,-7000.7,-353.40,-3074.4,-2951.7,-14030.,-1716.5,-1416.8,-5339.5,-3021.6,-5797.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
469.0000000000,5674.1,1112.8,1364.6,1640.7,1664.7,1201.7,2915.1,668.23,1650.9,358.67,607.47,769.16,0.0000,-4003.8,-6995.1,-352.66,-3073.1,-2948.9,-14028.,-1716.4,-1414.2,-5338.8,-3020.9,-5796.6,460.29,205.74,157.60,147.92,286.74,98.809,354.18,102.35,156.47,46.703,67.121,80.850,0.0000,-0.50703,-0.53574,-0.74516E-01,-0.46416,-0.38469,-1.8353,-1.4624,-0.14903,-1.3161,-0.17315,-1.8212
470.0000000000,5684.2,1113.7,1365.7,1642.6,1664.6,1202.8,2917.4,658.94,1645.9,357.95,606.14,763.72,0.0000,-3998.6,-6989.9,-352.04,-3071.8,-2946.2,-14027.,-1716.2,-1411.8,-5338.1,-3020.2,-5796.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
471.0000000000,5694.5,1115.2,1364.5,1652.5,1666.0,1191.6,2927.9,650.57,1644.7,358.24,607.57,754.77,0.0000,-3993.7,-6985.3,-351.51,-3070.5,-2943.6,-14025.,-1716.0,-1409.6,-5337.5,-3019.5,-5795.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
472.0000000000,5706.4,1106.4,1369.8,1619.3,1666.0,1161.4,2922.3,648.43,1648.8,357.73,595.67,744.33,0.0000,-3989.0,-6980.9,-351.03,-3069.2,-2941.1,-14023.,-1715.8,-1407.7,-5336.9,-3018.8,-5795.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
473.0000000000,5713.0,1104.4,1375.6,1625.7,1666.3,1160.7,2891.2,628.58,1660.9,357.01,592.25,743.15,0.0000,-3984.4,-6976.9,-350.60,-3067.9,-2938.6,-14022.,-1715.7,-1405.9,-5336.2,-3018.1,-5794.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
474.0000000000,5754.3,1100.2,1371.7,1593.1,1666.4,1163.0,2882.8,614.98,1622.0,357.72,588.98,743.68,0.0000,-3980.0,-6973.0,-350.20,-3066.6,-2936.1,-14020.,-1715.6,-1404.2,-5335.8,-3017.5,-5794.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
475.0000000000,5750.2,1108.2,1377.7,1591.7,1665.2,1178.0,2875.6,602.08,1625.6,357.11,586.86,743.07,0.0000,-4022.5,-6992.9,-353.97,-3065.7,-2961.8,-14019.,-1716.0,-1427.9,-5346.9,-3019.5,-5801.7,4005.4,1790.3,1371.4,1287.1,2495.2,859.83,3082.0,890.63,1361.6,406.41,584.08,703.55,0.0000,-4.4028,-4.6448,-0.64844,-4.0377,-3.3328,-15.956,-12.723,-1.2969,-11.450,-1.5043,-15.845
476.0000000000,5764.5,1103.9,1375.1,1590.0,1664.5,1164.8,2804.3,592.58,1626.1,356.47,586.06,743.85,0.0000,-3996.0,-6991.0,-353.37,-3064.5,-2942.2,-14018.,-1715.8,-1416.0,-5338.5,-3017.4,-5796.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
477.0000000000,5777.9,1094.3,1372.0,1592.4,1659.9,1151.4,2793.4,591.74,1629.2,355.90,585.43,742.71,0.0000,-3987.6,-6985.7,-352.29,-3063.3,-2937.5,-14016.,-1715.6,-1411.2,-5335.9,-3016.3,-5794.2,5.4394,2.4313,1.8624,1.7480,3.3885,1.1677,4.1854,1.2095,1.8490,0.55191,0.79319,0.95543,0.0000,-0.59707E-02,-0.63014E-02,-0.88058E-03,-0.54779E-02,-0.45115E-02,-0.21663E-01,-0.17277E-01,-0.17612E-02,-0.15548E-01,-0.20416E-02,-0.21516E-01
478.0000000000,5786.1,1098.5,1369.1,1605.3,1661.1,1146.0,2783.1,593.31,1628.5,355.31,575.79,734.86,0.0000,-3981.8,-6980.2,-351.35,-3062.1,-2934.4,-14014.,-1715.4,-1408.2,-5334.7,-3015.4,-5793.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
479.0000000000,5754.7,1096.5,1367.6,1609.7,1672.6,1130.4,2760.1,587.28,1589.9,354.82,564.55,735.28,0.0000,-3976.5,-6975.0,-350.59,-3060.8,-2931.5,-14013.,-1715.2,-1405.9,-5333.8,-3014.6,-5792.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
480.0000000000,5752.9,1089.5,1365.9,1610.2,1705.3,1127.3,2759.6,579.33,1585.6,353.48,562.49,731.76,0.0000,-3971.7,-6970.3,-349.96,-3059.6,-2928.9,-14011.,-1715.0,-1403.7,-5333.0,-3013.9,-5792.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
481.0000000000,5756.3,1101.4,1369.9,1603.8,1711.0,1129.4,2761.0,567.25,1582.4,353.33,563.28,731.39,0.0000,-3967.1,-6965.8,-349.43,-3058.3,-2926.3,-14009.,-1714.9,-1401.8,-5332.4,-3013.2,-5791.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
482.0000000000,5756.7,1100.6,1366.1,1619.2,1712.3,1133.8,2730.5,551.91,1576.8,354.00,562.91,728.73,0.0000,-3962.8,-6961.5,-348.96,-3057.1,-2923.8,-14007.,-1714.8,-1400.0,-5331.7,-3012.5,-5791.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
483.0000000000,5763.4,1099.7,1359.5,1616.2,1715.2,1138.9,2705.7,551.77,1544.0,353.66,562.30,723.69,0.0000,-3958.6,-6957.4,-348.55,-3055.8,-2921.4,-14006.,-1714.6,-1398.4,-5331.1,-3011.8,-5790.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
484.0000000000,5774.9,1098.9,1358.1,1585.0,1716.4,1142.2,2711.6,551.18,1542.8,353.62,560.03,715.24,0.0000,-3954.5,-6953.6,-348.16,-3054.6,-2919.0,-14004.,-1714.5,-1396.8,-5330.5,-3011.1,-5790.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
485.0000000000,5779.3,1080.8,1356.9,1587.0,1717.9,1141.1,2697.5,522.15,1545.0,352.26,551.24,710.20,0.0000,-3950.5,-6950.1,-347.81,-3053.4,-2916.6,-14002.,-1714.4,-1395.4,-5329.9,-3010.4,-5789.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
486.0000000000,5844.9,1076.4,1348.8,1586.9,1704.1,1140.0,2631.0,515.30,1546.8,350.45,549.24,710.33,0.0000,-3946.7,-6946.8,-347.46,-3052.2,-2914.3,-14000.,-1714.3,-1394.0,-5329.3,-3009.7,-5789.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
487.0000000000,5892.7,1086.7,1339.3,1587.8,1705.1,1139.7,2609.0,512.20,1544.1,350.35,548.18,707.17,0.0000,-3942.9,-6943.6,-347.13,-3051.0,-2912.0,-13999.,-1714.2,-1392.6,-5328.7,-3009.0,-5789.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
488.0000000000,5901.3,1087.3,1331.6,1589.1,1713.8,1140.6,2605.1,502.48,1540.8,349.26,542.75,701.41,0.0000,-3939.3,-6940.6,-346.81,-3049.8,-2909.8,-13997.,-1714.1,-1391.4,-5328.1,-3008.3,-5788.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
489.0000000000,5932.9,1096.0,1338.0,1589.2,1718.6,1138.0,2608.0,485.80,1546.7,348.32,537.90,703.23,0.0000,-3935.7,-6937.6,-346.48,-3048.7,-2907.6,-13996.,-1714.0,-1390.2,-5327.5,-3007.7,-5788.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
490.0000000000,5945.5,1089.7,1340.6,1589.5,1723.2,1137.1,2569.9,474.37,1550.0,345.02,538.75,702.92,0.0000,-3932.2,-6934.8,-346.16,-3047.7,-2905.4,-13994.,-1713.9,-1389.0,-5327.0,-3007.0,-5787.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
491.0000000000,5942.1,1088.8,1345.5,1590.7,1720.7,1140.3,2567.1,473.08,1549.7,342.29,540.98,703.53,0.0000,-3928.8,-6932.1,-345.84,-3046.8,-2903.2,-13993.,-1713.8,-1388.0,-5326.4,-3006.3,-5787.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
492.0000000000,5924.6,1096.0,1347.7,1594.7,1801.0,1131.4,2551.6,468.86,1548.5,343.86,541.01,706.39,0.0000,-3971.9,-6952.9,-349.66,-3046.2,-2929.1,-13992.,-1717.0,-1411.5,-5338.1,-3008.3,-5795.8,24033.,10742.,8228.9,7723.1,14971.,5159.1,18493.,5343.9,8169.5,2438.5,3504.6,4221.4,0.0000,-26.167,-27.551,-3.8907,-24.134,-19.626,-95.540,-76.307,-7.7814,-68.659,-8.9825,-95.010
493.0000000000,5911.1,1088.4,1338.0,1588.3,1834.2,1122.5,2546.9,462.86,1536.6,345.32,540.95,706.15,0.0000,-3946.4,-6952.0,-349.11,-3045.4,-2909.8,-13990.,-1716.1,-1400.6,-5329.9,-3006.2,-5790.6,0.63844,0.28537,0.21860,0.20517,0.39772,0.13705,0.49126,0.14196,0.21703,0.64779E-01,0.93099E-01,0.11214,0.0000,-0.69479E-03,-0.73175E-03,-0.10336E-03,-0.64081E-03,-0.52050E-03,-0.25378E-02,-0.20271E-02,-0.20672E-03,-0.18239E-02,-0.23855E-03,-0.25238E-02
494.0000000000,5921.0,1098.3,1354.0,1556.9,1832.3,1134.2,2553.6,454.64,1527.0,345.52,541.11,706.55,0.0000,-3985.6,-6971.1,-352.20,-3044.8,-2933.6,-13989.,-1716.9,-1421.4,-5339.2,-3007.8,-5797.1,11045.,4937.0,3781.9,3549.5,6880.8,2371.1,8499.0,2456.0,3754.6,1120.7,1610.7,1940.1,0.0000,-12.046,-12.667,-1.7881,-11.099,-9.0220,-43.900,-35.069,-3.5763,-31.553,-4.1263,-43.662
495.0000000000,5946.0,1100.2,1380.3,1531.7,1832.3,1121.4,2532.0,453.25,1532.1,342.28,541.08,705.91,0.0000,-4005.0,-6991.5,-355.19,-3044.4,-2941.6,-13987.,-1718.8,-1434.2,-5342.3,-3008.2,-5799.7,21147.,9452.1,7240.5,6795.5,13173.,4539.5,16272.,4702.1,7188.3,2145.6,3083.7,3714.4,0.0000,-23.115,-24.277,-3.4234,-21.271,-17.300,-84.037,-67.140,-6.8469,-60.407,-7.8984,-83.590
496.0000000000,5976.4,1105.1,1377.1,1509.5,1838.9,1081.3,2514.8,454.20,1532.0,337.32,533.86,696.38,0.0000,-3974.0,-6986.7,-353.45,-3043.7,-2919.7,-13985.,-1717.3,-1417.9,-5331.6,-3005.5,-5792.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
497.0000000000,5979.3,1086.2,1375.6,1480.7,1866.9,1076.4,2510.5,454.32,1530.5,338.47,532.40,692.85,0.0000,-3963.6,-6978.2,-351.49,-3042.7,-2914.1,-13983.,-1716.3,-1411.1,-5328.1,-3004.1,-5789.9,949.68,424.49,325.17,305.18,591.61,203.87,730.75,211.17,322.83,96.360,138.49,166.81,0.0000,-1.0366,-1.0897,-0.15375,-0.95397,-0.77390,-3.7732,-3.0151,-0.30749,-2.7127,-0.35448,-3.7537
498.0000000000,5976.7,1081.7,1380.8,1447.1,1871.7,1084.7,2506.4,441.51,1537.3,339.31,531.16,694.30,0.0000,-4003.2,-6993.3,-354.06,-3042.1,-2938.6,-13982.,-1718.5,-1432.3,-5338.5,-3005.8,-5797.1,23244.,10390.,7958.8,7469.6,14480.,4989.8,17886.,5168.5,7901.5,2358.5,3389.6,4082.9,0.0000,-25.422,-26.685,-3.7630,-23.374,-18.976,-92.341,-73.797,-7.5261,-66.393,-8.6743,-91.870
499.0000000000,5987.9,1081.3,1382.3,1421.3,1873.3,1089.7,2510.2,435.47,1545.4,337.94,531.49,683.89,0.0000,-4021.5,-7011.0,-356.75,-3041.6,-2946.5,-13981.,-1717.8,-1444.3,-5341.3,-3006.1,-5799.3,5336.3,2385.2,1827.1,1714.8,3324.3,1145.5,4106.1,1186.6,1814.0,541.44,778.15,937.32,0.0000,-5.8483,-6.1326,-0.86389,-5.3711,-4.3630,-21.196,-16.941,-1.7278,-15.242,-1.9910,-21.090
500.0000000000,5982.1,1078.9,1374.5,1423.6,1878.9,1082.2,2503.9,436.64,1543.8,335.92,531.98,680.95,0.0000,-3989.1,-7004.0,-354.82,-3040.7,-2924.3,-13979.,-1716.5,-1426.7,-5330.3,-3003.3,-5791.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
501.0000000000,5966.4,1077.8,1372.1,1423.8,1874.0,1085.1,2501.0,430.29,1545.3,334.58,533.03,679.22,0.0000,-3977.5,-6993.6,-352.72,-3039.7,-2918.5,-13977.,-1715.4,-1419.0,-5326.6,-3001.9,-5788.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
502.0000000000,5955.4,1082.2,1371.3,1420.6,1869.2,1077.2,2477.0,429.06,1532.3,332.54,526.37,679.65,0.0000,-3969.1,-6983.6,-351.03,-3038.6,-2914.6,-13975.,-1714.6,-1413.8,-5324.6,-3000.8,-5787.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
503.0000000000,5924.4,1083.4,1375.4,1419.0,1862.0,1073.6,2459.4,424.67,1528.5,331.99,519.72,668.27,0.0000,-3961.9,-6974.6,-349.72,-3037.5,-2911.2,-13973.,-1714.0,-1409.6,-5323.2,-2999.8,-5786.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
504.0000000000,5930.4,1096.6,1375.1,1421.2,1856.9,1075.0,2443.0,418.78,1529.5,332.72,516.93,671.10,0.0000,-3955.5,-6966.7,-348.70,-3036.4,-2908.1,-13972.,-1713.6,-1406.1,-5322.0,-2998.8,-5785.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
505.0000000000,5944.2,1096.9,1380.8,1423.0,1861.8,1046.4,2431.0,418.97,1532.1,326.46,512.13,677.41,0.0000,-3949.6,-6959.6,-347.86,-3035.2,-2905.2,-13970.,-1713.2,-1403.0,-5321.0,-2997.9,-5784.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
506.0000000000,5957.4,1098.9,1384.3,1423.5,1882.9,1040.8,2393.4,419.63,1542.4,322.80,496.02,679.90,0.0000,-3944.0,-6953.3,-347.16,-3034.2,-2902.5,-13968.,-1712.9,-1400.2,-5320.1,-2997.1,-5783.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
507.0000000000,5963.9,1103.7,1392.3,1428.1,1896.1,1042.7,2365.0,419.15,1554.1,321.68,494.30,670.44,0.0000,-3938.8,-6947.6,-346.56,-3033.2,-2900.0,-13967.,-1712.7,-1397.7,-5319.4,-2996.2,-5782.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
508.0000000000,5975.4,1111.9,1404.4,1443.1,1903.1,1058.6,2357.3,417.16,1545.2,321.01,492.74,670.08,0.0000,-3980.7,-6965.8,-350.16,-3032.5,-2925.5,-13966.,-1713.8,-1420.6,-5330.4,-2998.2,-5790.0,9177.8,4102.3,3142.5,2949.3,5717.3,1970.2,7062.0,2040.7,3119.8,931.22,1338.3,1612.1,0.0000,-10.007,-10.502,-1.4858,-9.2140,-7.4294,-36.425,-29.131,-2.9716,-26.205,-3.4148,-36.260
509.0000000000,5977.5,1111.9,1392.2,1435.0,1904.0,1052.3,2355.1,416.11,1526.6,315.68,492.68,669.54,0.0000,-3953.9,-6962.7,-349.44,-3031.7,-2905.9,-13964.,-1713.4,-1408.1,-5321.9,-2996.0,-5784.3,387.98,173.42,132.84,124.68,241.69,83.286,298.54,86.270,131.89,39.366,56.576,68.149,0.0000,-0.42279,-0.44386,-0.62810E-01,-0.38931,-0.31355,-1.5397,-1.2315,-0.12562,-1.1077,-0.14432,-1.5328
510.0000000000,5983.9,1122.0,1400.3,1443.5,1910.1,1031.3,2333.6,400.79,1538.9,311.24,493.71,658.97,0.0000,-3992.2,-6979.7,-352.39,-3031.1,-2929.3,-13963.,-1716.1,-1428.4,-5331.4,-2997.6,-5791.0,22822.,10201.,7814.3,7334.0,14217.,4899.2,17561.,5074.7,7758.0,2315.7,3328.0,4008.8,0.0000,-24.921,-26.124,-3.6947,-22.927,-18.480,-90.565,-72.441,-7.3894,-65.161,-8.4882,-90.166
511.0000000000,6002.2,1126.3,1403.0,1448.3,1912.2,1028.7,2333.2,398.47,1546.7,312.21,492.20,656.09,0.0000,-4010.6,-6998.5,-355.26,-3030.6,-2937.0,-13962.,-1735.6,-1440.3,-5338.3,-2997.9,-5798.6,0.15242E+06,68128.,52188.,48980.,94950.,32719.,0.11728E+06,33891.,51812.,15465.,22226.,26773.,0.0000,-166.79,-174.62,-24.675,-153.27,-123.62,-604.79,-483.88,-49.350,-435.17,-56.679,-602.18
512.0000000000,5988.2,1136.8,1411.2,1450.7,1911.1,1029.4,2335.2,397.95,1547.5,313.13,492.91,652.62,0.0000,-4025.6,-7015.8,-357.58,-3030.1,-2942.9,-13961.,-1731.0,-1449.5,-5341.1,-2997.9,-5802.0,9753.2,4359.5,3339.5,3134.2,6075.8,2093.7,7504.7,2168.7,3315.4,989.61,1422.2,1713.2,0.0000,-10.696,-11.185,-1.5789,-9.8155,-7.9210,-38.699,-30.965,-3.1579,-27.847,-3.6263,-38.536
513.0000000000,5991.3,1155.4,1427.4,1445.6,1920.5,1042.7,2329.1,399.36,1530.6,317.06,495.94,662.80,0.0000,-3992.5,-7007.6,-355.29,-3029.8,-2921.3,-13960.,-1725.8,-1430.4,-5329.8,-2995.5,-5794.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
514.0000000000,6001.4,1187.7,1440.9,1447.9,1924.5,1029.2,2345.6,392.85,1525.3,318.86,505.91,664.17,0.0000,-3982.1,-6997.6,-352.94,-3029.2,-2916.0,-13960.,-1721.8,-1421.9,-5325.5,-2994.9,-5790.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
515.0000000000,5998.2,1177.0,1428.3,1437.8,1927.4,1019.8,2341.3,380.85,1455.3,318.39,500.93,656.51,0.0000,-3973.7,-6987.4,-351.09,-3028.2,-2911.8,-13959.,-1718.8,-1416.2,-5323.6,-2994.2,-5787.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
516.0000000000,6040.6,1188.3,1433.5,1408.2,1930.0,1012.0,2335.7,378.15,1447.3,314.02,498.06,654.59,0.0000,-3966.4,-6977.4,-349.67,-3027.3,-2908.1,-13958.,-1716.7,-1411.5,-5321.6,-2993.4,-5785.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
517.0000000000,6080.9,1188.2,1429.0,1402.1,1932.6,957.84,2335.2,368.32,1440.8,310.88,501.86,652.50,0.0000,-3959.7,-6968.7,-348.55,-3026.4,-2904.5,-13956.,-1715.3,-1407.6,-5320.2,-2993.1,-5783.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
518.0000000000,6078.9,1186.0,1432.4,1399.2,1928.0,962.88,2314.8,365.78,1439.6,304.41,501.65,645.30,0.0000,-3953.4,-6960.1,-347.66,-3025.5,-2901.2,-13954.,-1714.2,-1404.1,-5318.9,-2992.5,-5781.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
519.0000000000,6093.6,1177.1,1430.7,1404.1,1919.6,929.46,2265.0,364.68,1442.0,301.36,499.84,640.55,0.0000,-3947.7,-6952.7,-346.93,-3024.6,-2898.2,-13952.,-1713.4,-1401.0,-5317.5,-2991.9,-5780.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
520.0000000000,6100.3,1169.4,1436.3,1406.1,1922.1,919.86,2266.8,362.58,1443.7,299.96,498.54,633.06,0.0000,-3942.2,-6946.2,-346.33,-3023.4,-2895.3,-13951.,-1712.9,-1398.3,-5316.5,-2991.5,-5779.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
521.0000000000,6105.8,1164.8,1437.4,1408.1,1915.5,916.19,2259.4,358.39,1445.3,298.26,490.82,628.77,0.0000,-3936.9,-6941.4,-345.82,-3022.1,-2892.5,-13950.,-1712.4,-1395.8,-5315.7,-2991.4,-5778.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
522.0000000000,6113.2,1163.9,1403.3,1401.4,1919.6,913.61,2267.6,358.51,1444.7,296.67,484.45,628.52,0.0000,-3931.9,-6936.5,-345.37,-3020.9,-2889.7,-13948.,-1712.1,-1393.5,-5315.0,-2991.3,-5777.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
523.0000000000,6156.4,1170.1,1391.9,1366.0,1928.3,913.86,2256.1,357.44,1453.9,294.86,484.47,629.62,0.0000,-3927.1,-6931.2,-344.94,-3019.7,-2887.1,-13947.,-1711.8,-1391.4,-5314.1,-2991.3,-5776.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
524.0000000000,6187.0,1169.3,1395.7,1362.2,1947.3,920.52,2249.2,355.20,1455.3,285.50,483.02,621.83,0.0000,-3922.5,-6927.1,-344.53,-3018.6,-2884.5,-13945.,-1711.6,-1389.4,-5313.1,-2991.0,-5775.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
525.0000000000,6185.3,1165.4,1404.3,1367.4,1937.0,922.74,2222.2,349.92,1467.2,283.59,479.29,624.00,0.0000,-3964.6,-6946.6,-348.26,-3017.9,-2910.0,-13945.,-1711.8,-1412.4,-5323.8,-2993.2,-5783.5,2236.8,999.82,765.89,718.81,1393.4,480.17,1721.2,497.37,760.36,226.96,326.18,392.90,0.0000,-2.4327,-2.5487,-0.36212,-2.2430,-1.7902,-8.8646,-7.1046,-0.72424,-6.3874,-0.82913,-8.8454
526.0000000000,6191.2,1175.9,1414.0,1372.2,1930.0,938.49,2212.7,344.41,1460.9,281.64,478.48,621.77,0.0000,-3985.2,-6967.5,-351.78,-3017.3,-2918.6,-13944.,-1711.8,-1426.1,-5326.6,-2993.5,-5785.8,1600.9,715.58,548.15,514.46,997.30,343.66,1231.9,355.98,544.20,162.44,233.45,281.20,0.0000,-1.7449,-1.8256,-0.25917,-1.6070,-1.2835,-6.3436,-5.0847,-0.51835,-4.5714,-0.59329,-6.3304
527.0000000000,6194.5,1167.0,1411.6,1370.9,1927.3,934.60,2206.6,342.12,1444.4,277.90,470.92,621.32,0.0000,-3954.6,-6963.1,-350.43,-3016.5,-2896.7,-13942.,-1711.6,-1410.5,-5315.9,-2990.9,-5778.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
528.0000000000,6196.8,1182.7,1427.7,1379.2,1921.2,945.18,2214.0,341.53,1447.9,270.13,463.38,619.81,0.0000,-3991.2,-6978.6,-352.85,-3015.9,-2919.2,-13941.,-1712.1,-1429.5,-5324.1,-2992.3,-5784.3,4867.7,2175.8,1666.7,1564.3,3032.4,1044.9,3745.6,1082.4,1654.7,493.91,709.83,855.03,0.0000,-5.3123,-5.5541,-0.78804,-4.8880,-3.9007,-19.283,-15.460,-1.5761,-13.899,-1.8029,-19.246
529.0000000000,6208.5,1188.5,1429.3,1384.2,1924.9,929.06,2214.5,331.09,1446.9,269.73,460.91,617.07,0.0000,-4008.5,-6995.6,-355.34,-3015.3,-2926.6,-13940.,-1715.9,-1440.7,-5327.0,-2992.5,-5787.1,30941.,13830.,10594.,9943.1,19275.,6642.1,23808.,6880.0,10518.,3139.5,4512.0,5434.9,0.0000,-33.835,-35.335,-5.0091,-31.097,-24.829,-122.56,-98.269,-10.018,-88.342,-11.457,-122.33
530.0000000000,6209.8,1189.4,1427.3,1388.1,1892.0,908.29,2222.2,328.36,1453.4,268.02,462.34,614.04,0.0000,-4022.6,-7011.4,-357.39,-3014.8,-2932.2,-13939.,-1722.4,-1449.2,-5329.5,-2992.4,-5790.2,57571.,25733.,19712.,18501.,35864.,12359.,44299.,12801.,19570.,5841.5,8395.3,10113.,0.0000,-63.081,-65.810,-9.3203,-57.905,-46.255,-228.00,-182.85,-18.641,-164.37,-21.313,-227.60
531.0000000000,6220.3,1185.3,1417.6,1386.8,1876.8,897.07,2224.1,327.82,1444.6,266.20,463.99,611.68,0.0000,-3988.4,-7001.8,-354.91,-3014.0,-2909.0,-13937.,-1719.4,-1429.7,-5318.7,-2989.5,-5783.3,654.95,292.75,224.25,210.47,408.01,140.60,503.96,145.63,222.64,66.455,95.507,115.04,0.0000,-0.71699,-0.74865,-0.10603,-0.65815,-0.52496,-2.5935,-2.0802,-0.21206,-1.8698,-0.24238,-2.5891
532.0000000000,6223.0,1183.4,1418.4,1383.4,1716.7,888.43,2225.8,327.15,1428.3,264.46,466.65,611.49,0.0000,-3975.6,-6989.0,-352.39,-3013.0,-2902.6,-13936.,-1716.9,-1420.7,-5314.7,-2987.9,-5780.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
533.0000000000,6225.2,1191.8,1410.9,1381.8,1688.1,881.44,2236.4,325.37,1429.2,263.15,468.50,610.55,0.0000,-3966.2,-6977.1,-350.42,-3011.8,-2898.2,-13935.,-1715.0,-1414.7,-5312.2,-2986.8,-5778.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
534.0000000000,6228.6,1198.7,1403.6,1377.6,1686.1,871.48,2248.4,318.76,1431.0,263.07,467.81,613.09,0.0000,-3958.2,-6966.5,-348.91,-3010.7,-2894.5,-13933.,-1713.6,-1409.8,-5310.4,-2985.7,-5776.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
535.0000000000,6228.9,1198.0,1400.3,1377.3,1690.7,883.90,2249.9,320.07,1435.3,263.86,467.13,613.52,0.0000,-3951.1,-6957.1,-347.74,-3009.6,-2891.4,-13932.,-1712.6,-1405.6,-5309.0,-2984.8,-5775.1,2.7208,1.2161,0.93160,0.87434,1.6949,0.58407,2.0936,0.60499,0.92488,0.27607,0.39676,0.47791,0.0000,-0.29656E-02,-0.31027E-02,-0.44047E-03,-0.27279E-02,-0.21667E-02,-0.10770E-01,-0.86410E-02,-0.88095E-03,-0.77666E-02,-0.10055E-02,-0.10755E-01
536.0000000000,6231.6,1207.2,1410.0,1380.5,1688.0,900.83,2257.2,321.63,1444.2,266.11,470.18,609.15,0.0000,-3991.7,-6972.2,-350.95,-3008.9,-2916.6,-13932.,-1757.1,-1427.6,-5328.8,-2986.8,-5793.9,0.33463E+06,0.14957E+06,0.11458E+06,0.10753E+06,0.20846E+06,71834.,0.25749E+06,74408.,0.11375E+06,33953.,48797.,58779.,0.0000,-365.47,-381.76,-54.174,-335.93,-267.09,-1324.5,-1063.2,-108.35,-955.24,-123.67,-1322.8
537.0000000000,6236.6,1314.0,1480.9,1383.7,1745.0,1000.9,2423.4,336.64,1434.7,289.96,504.20,655.25,0.0000,-4015.8,-6993.4,-354.18,-3010.1,-2930.0,-13937.,-1764.5,-1439.8,-5341.0,-2989.7,-5806.6,0.14116E+06,63097.,48334.,45363.,87939.,30303.,0.10862E+06,31389.,47986.,14323.,20585.,24796.,0.0000,-155.01,-161.37,-22.853,-142.12,-113.52,-559.78,-448.90,-45.706,-403.24,-52.277,-558.93
538.0000000000,6243.7,1373.3,1516.9,1379.1,1752.1,991.35,2438.3,348.94,1390.8,304.25,529.41,666.52,0.0000,-4037.2,-7015.7,-356.84,-3012.0,-2939.1,-13943.,-1756.6,-1448.9,-5350.2,-2994.1,-5811.4,46953.,20987.,16077.,15088.,29250.,10079.,36129.,10440.,15961.,4764.1,6846.8,8247.4,0.0000,-51.792,-53.762,-7.6013,-47.370,-37.953,-186.41,-149.42,-15.203,-134.21,-17.417,-186.17
539.0000000000,6251.2,1418.3,1482.0,1375.7,1769.4,934.98,2374.6,352.36,1398.1,300.45,548.82,687.22,0.0000,-4008.4,-7008.5,-354.85,-3013.9,-2916.6,-13945.,-1743.9,-1429.5,-5340.9,-2996.6,-5803.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
540.0000000000,6256.7,1424.2,1532.1,1349.6,1773.0,924.75,2309.3,361.72,1423.2,295.01,582.91,666.89,0.0000,-4044.7,-7023.3,-357.00,-3013.9,-2938.2,-13948.,-1734.8,-1447.6,-5347.2,-3004.3,-5805.8,2698.3,1206.1,923.91,867.12,1680.9,579.25,2076.3,599.99,917.25,273.79,393.48,473.97,0.0000,-2.9796,-3.0905,-0.43684,-2.7231,-2.1804,-10.712,-8.5923,-0.87367,-7.7165,-1.0013,-10.711
541.0000000000,6248.5,1442.4,1532.3,1345.8,1822.5,938.40,2265.1,367.90,1432.0,293.97,598.51,657.16,0.0000,-4061.7,-7040.0,-359.37,-3013.1,-2944.9,-13949.,-1744.3,-1457.7,-5349.6,-3010.6,-5808.8,0.12191E+06,54490.,41741.,39176.,75943.,26170.,93804.,27107.,41440.,12369.,17777.,21413.,0.0000,-134.84,-139.73,-19.736,-123.12,-98.600,-483.86,-388.29,-39.472,-348.66,-45.235,-484.06
542.0000000000,6278.5,1401.4,1519.1,1334.3,1785.9,926.74,2280.8,367.48,1421.8,291.16,568.14,653.29,0.0000,-4029.4,-7029.3,-357.22,-3011.7,-2921.0,-13949.,-1735.3,-1438.0,-5337.1,-3009.7,-5800.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
543.0000000000,6380.0,1421.5,1513.6,1321.9,1800.2,935.06,2385.8,360.47,1413.9,293.16,551.07,659.84,0.0000,-4019.1,-7014.9,-355.00,-3010.5,-2915.0,-13951.,-1728.5,-1428.9,-5331.0,-3008.4,-5795.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
544.0000000000,6368.6,1453.9,1559.4,1325.7,1809.3,938.09,2393.9,358.92,1411.1,299.26,544.44,655.15,0.0000,-4059.2,-7027.2,-357.42,-3009.5,-2938.5,-13955.,-1723.8,-1449.1,-5339.9,-3009.7,-5800.2,1655.1,739.79,566.70,531.86,1031.0,355.29,1273.5,368.02,562.61,167.93,241.35,290.72,0.0000,-1.8305,-1.8973,-0.26794,-1.6708,-1.3354,-6.5680,-5.2739,-0.53588,-4.7352,-0.61367,-6.5771
545.0000000000,6373.5,1433.4,1537.7,1325.7,1876.4,927.55,2307.4,356.58,1420.1,295.90,540.67,660.54,0.0000,-4030.6,-7017.8,-355.84,-3009.0,-2916.9,-13955.,-1720.3,-1432.6,-5329.5,-3007.1,-5792.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
546.0000000000,6381.1,1397.1,1530.5,1327.7,1899.4,914.59,2286.8,352.41,1421.8,293.14,542.70,645.20,0.0000,-4019.9,-7006.0,-354.10,-3008.1,-2910.4,-13956.,-1717.7,-1424.8,-5325.0,-3005.5,-5789.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
547.0000000000,6387.1,1397.9,1536.7,1329.8,1884.4,919.00,2277.8,362.67,1420.0,289.91,544.69,646.11,0.0000,-4010.8,-6995.0,-352.68,-3007.2,-2905.8,-13956.,-1715.9,-1419.3,-5322.6,-3005.4,-5787.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
548.0000000000,6387.8,1376.6,1533.0,1331.0,1877.7,910.62,2272.1,359.41,1412.9,278.95,537.65,654.60,0.0000,-4003.4,-6984.5,-351.54,-3006.5,-2901.7,-13955.,-1714.6,-1414.7,-5320.3,-3005.5,-5786.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
549.0000000000,6389.7,1350.6,1547.6,1333.1,1857.5,890.26,2340.1,358.69,1425.9,277.30,530.70,656.06,0.0000,-3996.4,-6975.5,-350.63,-3005.9,-2898.0,-13955.,-1713.7,-1410.7,-5319.3,-3004.6,-5785.5,316.52,141.48,108.38,101.72,197.18,67.947,243.56,70.381,107.60,32.116,46.157,55.598,0.0000,-0.34789,-0.36193,-0.51242E-01,-0.31853,-0.25305,-1.2546,-1.0086,-0.10248,-0.90551,-0.11709,-1.2576
550.0000000000,6388.5,1349.6,1568.1,1335.2,1859.0,880.44,2308.5,359.58,1412.0,282.03,523.26,663.04,0.0000,-3989.8,-6968.7,-349.88,-3005.2,-2894.6,-13955.,-1713.0,-1407.8,-5318.7,-3003.5,-5785.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
551.0000000000,6387.0,1353.2,1569.8,1334.9,1912.3,884.12,2279.4,360.56,1420.7,278.96,523.68,652.08,0.0000,-3984.5,-6962.6,-349.23,-3004.8,-2891.5,-13955.,-1712.5,-1405.3,-5317.6,-3002.4,-5784.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
552.0000000000,6376.7,1344.8,1573.1,1341.3,1893.6,879.21,2295.4,360.21,1406.4,265.85,531.22,644.48,0.0000,-3979.1,-6956.2,-348.63,-3005.0,-2888.8,-13955.,-1712.2,-1402.7,-5317.2,-3002.0,-5784.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
553.0000000000,6358.2,1347.1,1583.7,1346.1,1887.7,897.42,2320.7,356.25,1415.6,268.44,519.74,645.21,0.0000,-3974.0,-6950.9,-348.06,-3005.7,-2886.1,-13954.,-1711.9,-1400.5,-5317.6,-3000.7,-5783.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
554.0000000000,6351.0,1358.1,1579.1,1349.1,1903.7,909.44,2317.9,343.23,1442.9,267.28,513.47,629.48,0.0000,-3969.9,-6945.1,-347.53,-3006.7,-2883.5,-13954.,-1711.6,-1398.4,-5317.5,-2998.6,-5782.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
555.0000000000,6381.0,1378.9,1562.6,1346.6,1884.0,912.36,2314.1,340.20,1457.0,266.33,506.24,625.44,0.0000,-3965.9,-6939.7,-347.04,-3007.4,-2880.8,-13954.,-1711.4,-1395.8,-5317.3,-2996.6,-5781.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
556.0000000000,6393.6,1386.8,1585.9,1304.2,1867.1,928.69,2287.6,338.77,1444.1,260.83,497.95,623.65,0.0000,-4008.7,-6961.1,-350.70,-3007.6,-2906.2,-13954.,-1711.5,-1418.5,-5327.3,-2997.6,-5789.2,1484.8,663.67,508.39,477.14,924.95,318.73,1142.5,330.15,504.72,150.65,216.51,260.80,0.0000,-1.6264,-1.6929,-0.24037,-1.4932,-1.1821,-5.8813,-4.7294,-0.48074,-4.2460,-0.54796,-5.8948
557.0000000000,6398.6,1353.5,1573.4,1313.0,1900.4,936.94,2263.9,341.70,1426.5,259.19,504.22,621.59,0.0000,-4028.7,-6982.7,-354.14,-3009.5,-2915.8,-13954.,-1711.7,-1431.9,-5330.1,-2997.7,-5791.6,1825.8,816.10,625.15,586.73,1137.4,391.94,1404.9,405.98,620.64,185.25,266.24,320.70,0.0000,-2.0042,-2.0835,-0.29558,-1.8381,-1.4567,-7.2311,-5.8152,-0.59116,-5.2209,-0.67364,-7.2477
558.0000000000,6410.7,1349.3,1594.4,1313.1,1902.2,922.46,2233.0,337.58,1419.3,263.24,514.13,622.23,0.0000,-4044.6,-7001.2,-356.87,-3010.5,-2922.3,-13953.,-1714.9,-1441.9,-5331.9,-2998.2,-5793.4,25347.,11330.,8678.7,8145.3,15790.,5441.1,19504.,5636.0,8616.1,2571.8,3696.2,4452.2,0.0000,-27.881,-28.954,-4.1034,-25.542,-20.259,-100.37,-80.727,-8.2068,-72.474,-9.3499,-100.60
559.0000000000,6427.7,1348.4,1577.7,1307.2,1879.4,895.10,2217.6,333.73,1399.5,257.28,506.88,617.99,0.0000,-4011.4,-6993.8,-354.85,-3011.0,-2899.7,-13952.,-1713.9,-1424.0,-5320.8,-2995.7,-5786.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
560.0000000000,6483.1,1334.5,1572.0,1304.0,1889.9,892.73,2220.0,333.32,1393.8,255.28,510.18,615.83,0.0000,-3999.2,-6982.7,-352.66,-3011.2,-2893.8,-13950.,-1713.0,-1416.1,-5317.1,-2994.5,-5783.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
561.0000000000,6543.7,1351.0,1568.2,1297.8,1878.7,886.28,2233.7,335.38,1390.6,254.25,503.76,614.37,0.0000,-3990.3,-6972.0,-350.90,-3011.1,-2889.9,-13949.,-1712.3,-1410.8,-5315.0,-2993.6,-5781.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
562.0000000000,6362.0,1374.1,1565.3,1306.8,1868.2,901.47,2210.3,339.40,1391.1,254.63,501.44,613.53,0.0000,-4029.8,-6986.1,-353.69,-3011.3,-2914.8,-13949.,-1716.3,-1432.5,-5326.0,-2995.5,-5789.8,33237.,14856.,11380.,10681.,20705.,7134.9,25575.,7390.5,11298.,3372.4,4846.7,5838.1,0.0000,-36.523,-37.946,-5.3808,-33.470,-26.494,-131.56,-105.83,-10.762,-95.005,-12.247,-131.85
563.0000000000,6338.0,1368.2,1550.3,1316.0,1879.9,899.69,2190.1,337.19,1394.4,255.77,503.19,612.03,0.0000,-4047.9,-7003.1,-356.53,-3011.6,-2922.9,-13949.,-1720.3,-1444.6,-5330.1,-2995.5,-5793.7,39916.,17842.,13667.,12827.,24866.,8568.7,30714.,8875.6,13569.,4050.1,5820.7,7011.3,0.0000,-43.949,-45.606,-6.4620,-40.236,-31.876,-157.99,-127.10,-12.924,-114.09,-14.706,-158.32
564.0000000000,6341.8,1373.6,1548.7,1300.3,1876.8,906.41,2172.2,335.54,1410.2,253.77,506.02,608.33,0.0000,-4062.4,-7018.6,-358.84,-3011.9,-2928.9,-13949.,-1721.8,-1453.5,-5332.0,-2995.0,-5795.9,29627.,13242.,10144.,9520.6,18456.,6359.9,22797.,6587.7,10071.,3006.1,4320.2,5204.0,0.0000,-32.685,-33.880,-4.7963,-29.889,-23.697,-117.25,-94.333,-9.5925,-84.674,-10.914,-117.50
565.0000000000,6348.0,1361.7,1528.5,1292.5,1864.7,898.54,2165.0,335.22,1395.6,248.64,504.03,601.27,0.0000,-4027.8,-7008.1,-356.53,-3011.8,-2905.9,-13948.,-1718.8,-1434.0,-5320.3,-2991.6,-5788.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
566.0000000000,6353.1,1365.8,1531.5,1291.7,1837.0,899.55,2177.4,336.59,1387.2,246.73,505.62,601.95,0.0000,-4014.5,-6994.7,-354.13,-3011.5,-2899.8,-13948.,-1716.4,-1424.7,-5315.8,-2989.7,-5784.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
567.0000000000,6375.8,1376.4,1532.4,1290.1,1823.4,895.72,2184.3,339.19,1386.7,247.96,503.28,605.13,0.0000,-4004.3,-6982.0,-352.23,-3011.1,-2895.6,-13947.,-1714.6,-1418.5,-5313.3,-2988.4,-5782.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
568.0000000000,6373.4,1379.4,1534.2,1294.1,1820.6,898.70,2199.0,337.52,1361.3,248.90,506.72,602.19,0.0000,-3995.7,-6971.7,-350.77,-3010.3,-2892.5,-13946.,-1713.4,-1413.5,-5311.0,-2987.4,-5780.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
569.0000000000,6378.8,1386.8,1541.2,1298.5,1833.8,890.85,2202.6,328.35,1315.4,248.64,515.70,603.95,0.0000,-3988.7,-6963.5,-349.65,-3009.6,-2889.5,-13946.,-1712.4,-1409.3,-5309.4,-2986.9,-5778.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
570.0000000000,6436.2,1380.8,1540.8,1302.3,1848.8,886.33,2202.2,329.66,1289.1,249.04,515.12,605.34,0.0000,-3981.5,-6956.5,-348.77,-3008.9,-2886.4,-13946.,-1711.8,-1405.6,-5308.2,-2986.1,-5777.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
571.0000000000,6475.9,1383.4,1539.9,1313.2,1848.2,892.44,2204.2,335.02,1299.0,250.11,517.21,607.58,0.0000,-4021.6,-6972.5,-352.19,-3008.5,-2911.5,-13946.,-1713.3,-1427.8,-5319.4,-2988.3,-5785.2,14115.,6309.3,4833.1,4536.0,8793.2,3030.1,10861.,3138.6,4798.2,1432.2,2058.3,2479.4,0.0000,-15.506,-16.100,-2.2851,-14.216,-11.228,-55.850,-44.937,-4.5703,-40.331,-5.1950,-55.966
572.0000000000,6489.1,1370.5,1534.4,1324.7,1825.3,879.85,2177.7,336.35,1288.3,251.73,511.41,613.87,0.0000,-3992.5,-6967.1,-351.33,-3007.4,-2890.8,-13945.,-1712.4,-1414.2,-5311.3,-2986.0,-5779.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
573.0000000000,6494.5,1356.8,1529.0,1328.6,1823.7,835.59,2170.9,338.15,1289.3,249.73,503.58,617.23,0.0000,-3981.8,-6958.4,-350.04,-3006.3,-2885.2,-13944.,-1711.8,-1408.0,-5308.7,-2984.6,-5777.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
574.0000000000,6488.1,1347.3,1541.4,1335.1,1838.7,830.57,2172.4,338.58,1278.2,250.81,504.47,615.43,0.0000,-3973.8,-6949.9,-348.93,-3005.4,-2881.3,-13942.,-1711.3,-1403.8,-5307.2,-2983.2,-5776.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
575.0000000000,6491.1,1340.2,1543.1,1332.7,1829.6,825.46,2176.4,335.23,1235.8,251.31,503.18,615.54,0.0000,-3966.8,-6942.3,-348.03,-3004.6,-2877.8,-13941.,-1710.8,-1400.4,-5306.3,-2982.4,-5775.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
576.0000000000,6488.1,1321.3,1546.2,1338.9,1803.9,827.72,2156.7,333.47,1231.5,250.06,498.65,613.33,0.0000,-3960.1,-6935.5,-347.29,-3003.8,-2874.6,-13939.,-1710.5,-1397.3,-5305.6,-2981.5,-5774.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
577.0000000000,6473.0,1314.3,1558.3,1344.0,1807.4,819.35,2158.8,333.69,1236.8,249.57,490.37,611.77,0.0000,-3953.8,-6929.3,-346.66,-3002.8,-2871.3,-13938.,-1710.3,-1394.4,-5304.8,-2980.5,-5773.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
578.0000000000,6456.3,1313.3,1558.3,1342.2,1799.2,813.74,2163.2,331.55,1259.2,250.53,484.48,617.62,0.0000,-3947.7,-6923.6,-346.11,-3001.8,-2868.2,-13936.,-1710.1,-1391.8,-5304.3,-2979.6,-5772.8,78.904,35.268,27.017,25.356,49.154,16.938,60.714,17.545,26.822,8.0060,11.506,13.860,0.0000,-0.86011E-01,-0.89642E-01,-0.12774E-01,-0.79196E-01,-0.62146E-01,-0.31192,-0.25112,-0.25548E-01,-0.22537,-0.29012E-01,-0.31265
579.0000000000,6454.8,1323.6,1553.4,1346.7,1788.4,822.63,2175.7,328.15,1259.5,253.38,481.28,618.96,0.0000,-3988.5,-6941.7,-349.75,-3001.1,-2893.3,-13935.,-1717.9,-1414.3,-5317.0,-2981.4,-5782.2,59344.,26526.,20319.,19070.,36969.,12739.,45664.,13196.,20173.,6021.4,8653.8,10424.,0.0000,-64.802,-67.446,-9.6073,-59.634,-46.846,-234.56,-188.87,-19.215,-169.50,-21.820,-235.12
580.0000000000,6450.1,1341.9,1550.7,1359.1,1796.4,827.76,2174.4,328.43,1276.0,252.71,476.89,623.61,0.0000,-4007.5,-6961.6,-353.20,-3000.6,-2901.4,-13933.,-1736.8,-1427.4,-5325.2,-2981.8,-5791.1,0.15512E+06,69336.,53113.,49848.,96633.,33299.,0.11936E+06,34492.,52730.,15739.,22620.,27247.,0.0000,-169.72,-176.44,-25.112,-156.03,-122.68,-613.04,-493.75,-50.225,-443.03,-57.033,-614.55
581.0000000000,6434.7,1350.1,1527.6,1339.3,1788.5,827.45,2196.9,330.59,1272.6,252.63,471.94,631.67,0.0000,-3975.4,-6955.2,-351.79,-2999.7,-2879.2,-13932.,-1729.9,-1411.3,-5316.7,-2979.3,-5786.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
582.0000000000,6416.1,1384.6,1545.8,1326.1,1810.7,876.81,2269.6,333.51,1280.6,258.93,483.32,641.23,0.0000,-3965.8,-6945.8,-350.08,-2999.5,-2875.8,-13932.,-1724.3,-1404.2,-5313.3,-2979.0,-5784.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
583.0000000000,6424.3,1371.2,1560.9,1303.0,1804.0,852.59,2261.1,328.85,1288.0,257.68,484.86,632.10,0.0000,-3959.1,-6939.4,-348.69,-2998.7,-2872.4,-13935.,-1720.0,-1399.7,-5311.2,-2979.0,-5781.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
584.0000000000,6432.5,1375.7,1557.9,1298.1,1797.4,867.12,2224.0,329.63,1279.1,253.65,481.63,626.88,0.0000,-3952.8,-6931.8,-347.61,-2997.8,-2869.0,-13936.,-1716.9,-1396.1,-5309.5,-2978.8,-5779.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
585.0000000000,6446.5,1382.1,1545.6,1298.1,1887.2,862.26,2200.3,330.74,1288.2,254.04,483.27,624.96,0.0000,-3946.4,-6924.5,-346.72,-2996.9,-2865.2,-13936.,-1714.7,-1393.2,-5308.2,-2978.9,-5777.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
586.0000000000,6478.1,1395.6,1535.6,1297.1,1909.4,858.86,2211.6,330.86,1293.7,253.71,477.17,628.68,0.0000,-3940.3,-6917.2,-345.99,-2996.0,-2862.0,-13935.,-1713.2,-1391.0,-5306.6,-2978.7,-5775.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
587.0000000000,6478.5,1416.2,1547.5,1296.8,1917.3,865.84,2231.5,330.30,1282.2,253.79,492.20,620.98,0.0000,-3934.6,-6911.7,-345.40,-2994.7,-2859.1,-13934.,-1712.1,-1389.1,-5305.3,-2979.3,-5774.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
588.0000000000,6496.1,1431.0,1553.5,1300.0,1915.1,873.54,2225.6,335.13,1282.5,252.92,497.55,617.73,0.0000,-3929.1,-6907.3,-344.90,-2993.3,-2856.5,-13934.,-1711.3,-1387.4,-5304.2,-2979.8,-5773.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
589.0000000000,6492.0,1436.4,1544.5,1295.7,1913.9,899.50,2221.5,337.52,1279.4,252.01,508.60,619.20,0.0000,-3970.5,-6927.2,-348.57,-2992.3,-2882.1,-13934.,-1713.0,-1410.5,-5315.3,-2983.4,-5780.8,15980.,7142.7,5471.5,5135.2,9954.8,3430.4,12296.,3553.2,5432.0,1621.4,2330.2,2806.9,0.0000,-17.408,-18.110,-2.5870,-16.035,-12.554,-63.150,-50.882,-5.1740,-45.650,-5.8725,-63.356
590.0000000000,6494.6,1431.0,1532.5,1303.5,1897.7,915.69,2185.9,335.42,1280.1,252.23,500.60,620.88,0.0000,-3990.4,-6948.2,-352.03,-2991.5,-2890.6,-13933.,-1717.2,-1424.3,-5319.1,-2985.0,-5784.4,37517.,16770.,12846.,12056.,23372.,8053.7,28868.,8342.2,12753.,3806.7,5470.9,6590.0,0.0000,-40.956,-42.552,-6.0737,-37.684,-29.529,-148.25,-119.46,-12.147,-107.17,-13.785,-148.74
591.0000000000,6513.0,1399.5,1560.4,1303.0,1875.6,915.35,2164.3,333.31,1278.2,251.56,492.51,620.53,0.0000,-3959.8,-6943.6,-350.61,-2990.6,-2868.3,-13931.,-1715.2,-1408.8,-5308.6,-2982.2,-5777.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
592.0000000000,6541.6,1386.9,1558.1,1316.8,1864.4,885.49,2176.5,330.67,1274.0,247.30,486.20,622.78,0.0000,-3949.1,-6934.4,-348.82,-2989.4,-2862.2,-13929.,-1713.6,-1402.2,-5304.7,-2980.1,-5775.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
593.0000000000,6531.7,1371.8,1557.4,1332.8,1874.7,870.71,2187.6,323.47,1274.3,242.58,483.06,622.75,0.0000,-3941.1,-6925.4,-347.34,-2988.1,-2858.1,-13927.,-1712.3,-1397.7,-5302.6,-2978.5,-5773.5,1.7914,0.80073,0.61338,0.57568,1.1160,0.38456,1.3784,0.39833,0.60896,0.18177,0.26123,0.31467,0.0000,-0.19497E-02,-0.20294E-02,-0.29001E-03,-0.17953E-02,-0.14013E-02,-0.70755E-02,-0.57034E-02,-0.58003E-03,-0.51165E-02,-0.65745E-03,-0.70997E-02
594.0000000000,6522.2,1358.6,1565.8,1357.8,1874.4,876.39,2160.1,319.88,1279.3,243.04,480.46,627.81,0.0000,-3980.4,-6940.7,-350.31,-2987.2,-2882.8,-13927.,-1712.7,-1419.3,-5312.8,-2980.0,-5780.6,9429.2,4214.7,3228.6,3030.1,5874.0,2024.1,7255.5,2096.7,3205.3,956.74,1375.0,1656.3,0.0000,-10.279,-10.686,-1.5265,-9.4594,-7.3897,-37.236,-30.019,-3.0530,-26.929,-3.4596,-37.365
595.0000000000,6520.4,1382.2,1561.7,1370.0,1892.8,872.16,2142.8,320.49,1286.4,241.08,481.36,625.20,0.0000,-3998.5,-6958.0,-353.27,-2986.8,-2890.7,-13926.,-1718.2,-1431.6,-5316.7,-2980.3,-5784.2,47397.,21186.,16229.,15231.,29526.,10175.,36470.,10539.,16112.,4809.1,6911.6,8325.4,0.0000,-51.765,-53.756,-7.6731,-47.589,-37.203,-187.15,-150.89,-15.346,-135.36,-17.386,-187.80
596.0000000000,6511.9,1399.3,1570.1,1379.1,1908.6,866.49,2141.2,320.22,1292.1,240.86,486.21,623.00,0.0000,-4013.0,-6974.4,-355.66,-2986.9,-2896.6,-13924.,-1723.8,-1441.0,-5319.6,-2980.2,-5787.5,58663.,26221.,20086.,18851.,36544.,12593.,45139.,13044.,19941.,5952.2,8554.4,10304.,0.0000,-64.192,-66.595,-9.4969,-58.943,-46.108,-231.60,-186.76,-18.994,-167.52,-21.514,-232.41
597.0000000000,6501.4,1410.7,1557.6,1368.2,1905.4,843.77,2149.1,325.18,1276.0,238.70,490.92,623.14,0.0000,-3978.9,-6965.6,-353.39,-2986.7,-2873.6,-13923.,-1720.0,-1422.5,-5308.7,-2977.3,-5780.4,214.85,96.034,73.565,69.043,133.84,46.121,165.32,47.773,73.034,21.800,31.330,37.739,0.0000,-0.23488,-0.24389,-0.34782E-01,-0.21568,-0.16847,-0.84813,-0.68397,-0.69565E-01,-0.61349,-0.78769E-01,-0.85115
598.0000000000,6484.9,1423.0,1555.3,1345.4,1897.5,844.41,2180.1,326.97,1277.8,240.60,500.98,628.84,0.0000,-3966.3,-6953.7,-351.00,-2986.2,-2867.4,-13921.,-1716.9,-1414.2,-5304.5,-2975.9,-5777.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
599.0000000000,6495.6,1439.8,1550.6,1334.8,1906.2,873.10,2218.8,328.66,1263.4,243.52,508.06,634.46,0.0000,-3957.9,-6942.6,-349.11,-2986.0,-2864.3,-13921.,-1714.6,-1408.6,-5302.1,-2975.4,-5774.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
600.0000000000,6484.8,1432.0,1563.3,1333.4,1900.2,879.16,2219.3,327.14,1257.6,242.70,505.73,635.74,0.0000,-3950.9,-6933.9,-347.66,-2984.8,-2860.9,-13921.,-1712.9,-1404.1,-5300.3,-2974.7,-5773.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
601.0000000000,6493.2,1421.7,1564.0,1327.1,1932.0,879.15,2237.1,321.48,1251.5,243.08,498.37,632.08,0.0000,-3943.9,-6925.8,-346.52,-2983.5,-2857.6,-13920.,-1711.7,-1400.2,-5299.0,-2974.1,-5771.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
602.0000000000,6601.7,1416.8,1565.8,1330.6,1944.5,875.49,2223.5,319.08,1249.9,241.06,494.39,636.90,0.0000,-3937.3,-6918.1,-345.58,-2982.2,-2854.2,-13919.,-1710.9,-1396.7,-5297.9,-2973.4,-5770.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
603.0000000000,6595.7,1411.1,1568.7,1324.5,1948.7,880.56,2240.5,322.08,1249.3,239.60,493.48,636.30,0.0000,-3930.9,-6911.2,-344.80,-2981.1,-2850.8,-13918.,-1710.2,-1393.6,-5296.8,-2972.5,-5768.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
604.0000000000,6607.0,1397.0,1565.1,1324.2,1959.2,872.68,2213.6,324.22,1239.8,240.71,499.66,634.56,0.0000,-3925.0,-6904.5,-344.10,-2980.3,-2847.6,-13917.,-1709.8,-1390.8,-5296.3,-2972.0,-5767.8,2.6023,1.1632,0.89104,0.83627,1.6211,0.55864,2.0024,0.57865,0.88461,0.26405,0.37948,0.45710,0.0000,-0.28255E-02,-0.29420E-02,-0.42129E-03,-0.26032E-02,-0.20226E-02,-0.10273E-01,-0.82845E-02,-0.84259E-03,-0.74303E-02,-0.95251E-03,-0.10310E-01
605.0000000000,6611.9,1393.4,1561.1,1329.1,1969.7,867.60,2208.5,327.37,1227.0,239.83,499.70,635.62,0.0000,-3919.3,-6898.6,-343.49,-2979.4,-2844.6,-13915.,-1709.6,-1388.2,-5295.8,-2971.2,-5767.1,1225.5,547.77,419.61,393.82,763.43,263.07,942.97,272.50,416.58,124.34,178.70,215.26,0.0000,-1.3292,-1.3845,-0.19840,-1.2254,-0.95117,-4.8375,-3.9012,-0.39679,-3.4989,-0.44846,-4.8548
606.0000000000,6623.3,1399.7,1569.0,1326.4,1981.7,882.09,2216.6,333.62,1229.6,238.83,500.87,633.80,0.0000,-3913.7,-6894.5,-342.92,-2978.3,-2841.9,-13914.,-1709.3,-1385.9,-5294.9,-2970.6,-5766.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
607.0000000000,6629.2,1414.6,1577.8,1333.1,1964.6,894.97,2234.4,332.39,1232.7,236.00,497.49,636.55,0.0000,-3955.0,-6912.6,-346.50,-2977.6,-2867.4,-13914.,-1710.0,-1408.3,-5305.6,-2972.6,-5773.9,7172.3,3205.9,2455.8,2304.8,4468.0,1539.7,5518.9,1594.8,2438.1,727.74,1045.9,1259.8,0.0000,-7.7866,-8.1007,-1.1611,-7.1775,-5.5725,-28.307,-22.830,-2.3223,-20.476,-2.6237,-28.408
608.0000000000,6645.3,1408.9,1582.9,1335.0,1959.4,902.16,2246.5,327.82,1236.0,236.57,501.98,637.59,0.0000,-3974.4,-6932.9,-349.91,-2977.0,-2875.7,-13914.,-1709.9,-1421.7,-5308.5,-2973.4,-5776.1,1923.0,859.55,658.44,617.97,1198.0,412.81,1479.7,427.60,653.69,195.12,280.42,337.78,0.0000,-2.0920,-2.1737,-0.31132,-1.9262,-1.4967,-7.5886,-6.1209,-0.62264,-5.4897,-0.70337,-7.6158
609.0000000000,6677.7,1385.4,1580.8,1336.4,1944.4,891.39,2267.8,328.88,1224.3,237.91,503.36,636.97,0.0000,-3943.0,-6928.7,-348.45,-2976.2,-2853.7,-13912.,-1709.5,-1406.0,-5297.9,-2971.0,-5768.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
610.0000000000,6730.6,1385.7,1573.1,1335.5,1895.0,875.77,2274.1,328.83,1231.6,237.81,499.50,638.01,0.0000,-3931.9,-6920.0,-346.64,-2975.2,-2848.0,-13911.,-1709.2,-1399.2,-5294.7,-2969.7,-5766.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
611.0000000000,6790.4,1388.6,1573.4,1333.4,1890.5,868.28,2280.2,331.08,1231.4,239.20,501.03,642.25,0.0000,-3923.8,-6911.5,-345.12,-2974.2,-2844.2,-13910.,-1708.9,-1394.6,-5293.2,-2968.6,-5765.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
612.0000000000,6787.2,1373.6,1573.2,1329.7,1874.7,865.68,2283.5,335.46,1239.1,238.77,498.77,642.65,0.0000,-3916.8,-6903.5,-343.92,-2973.2,-2841.0,-13909.,-1708.7,-1391.0,-5292.2,-2967.7,-5764.1,882.84,394.61,302.28,283.70,549.97,189.52,679.32,196.31,300.11,89.578,128.74,155.07,0.0000,-0.95655,-0.99615,-0.14292,-0.88198,-0.68230,-3.4823,-2.8094,-0.28585,-2.5196,-0.32249,-3.4944
613.0000000000,6780.1,1370.5,1580.6,1340.3,1876.6,877.05,2286.2,338.30,1248.0,236.30,497.38,644.40,0.0000,-3957.0,-6920.2,-347.07,-2972.5,-2866.1,-13908.,-1714.9,-1413.0,-5304.1,-2969.5,-5773.0,47210.,21102.,16165.,15171.,29410.,10134.,36326.,10497.,16048.,4790.1,6884.3,8292.5,0.0000,-51.245,-53.291,-7.6428,-47.216,-36.568,-186.20,-150.23,-15.286,-134.73,-17.243,-186.84
614.0000000000,6790.1,1373.6,1579.3,1328.4,1882.9,881.97,2293.6,339.69,1249.5,235.71,500.69,645.46,0.0000,-3975.3,-6939.4,-350.16,-2972.1,-2874.4,-13908.,-1715.0,-1425.7,-5308.0,-2970.1,-5776.5,13294.,5942.1,4551.8,4272.1,8281.5,2853.8,10229.,2956.0,4519.0,1348.9,1938.6,2335.1,0.0000,-14.459,-15.018,-2.1522,-13.308,-10.316,-52.428,-42.302,-4.3043,-37.936,-4.8548,-52.608
615.0000000000,6794.7,1375.6,1567.5,1318.3,1870.3,870.53,2283.9,337.50,1239.0,235.75,499.48,645.79,0.0000,-3943.4,-6933.6,-348.48,-2971.3,-2852.2,-13906.,-1713.2,-1409.3,-5297.5,-2967.7,-5769.5,249.91,111.70,85.568,80.308,155.68,53.647,192.29,55.569,84.951,25.357,36.442,43.896,0.0000,-0.27159,-0.28230,-0.40458E-01,-0.24997,-0.19353,-0.98550,-0.79517,-0.80915E-01,-0.71310,-0.91237E-01,-0.98883
616.0000000000,6778.5,1385.9,1574.6,1322.5,1874.9,883.63,2273.8,335.19,1249.9,235.60,498.84,645.99,0.0000,-3978.9,-6947.7,-350.65,-2970.6,-2874.6,-13906.,-1716.4,-1427.6,-5306.4,-2969.1,-5775.9,35092.,15686.,12016.,11277.,21861.,7533.2,27002.,7803.0,11929.,3560.7,5117.3,6164.0,0.0000,-38.207,-39.665,-5.6811,-35.134,-27.227,-138.38,-111.66,-11.362,-100.13,-12.810,-138.84
617.0000000000,6612.7,1385.0,1571.7,1322.7,1868.2,872.86,2265.7,337.33,1249.9,235.07,500.94,645.53,0.0000,-3948.2,-6940.1,-348.79,-2969.5,-2853.6,-13905.,-1714.1,-1412.0,-5296.9,-2966.6,-5769.7,128.69,57.520,44.062,41.354,80.166,27.625,99.020,28.614,43.745,13.057,18.765,22.604,0.0000,-0.13998,-0.14543,-0.20833E-01,-0.12873,-0.99642E-01,-0.50742,-0.40944,-0.41666E-01,-0.36716,-0.46960E-01,-0.50908
618.0000000000,6618.1,1383.9,1572.6,1324.4,1878.7,866.83,2262.2,337.42,1238.2,236.27,505.07,642.85,0.0000,-3936.6,-6929.8,-346.77,-2968.5,-2848.0,-13904.,-1712.3,-1404.7,-5293.5,-2965.4,-5766.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
619.0000000000,6620.8,1384.9,1575.5,1329.2,1880.3,863.36,2251.1,337.19,1228.6,236.35,504.80,639.22,0.0000,-3928.1,-6920.0,-345.11,-2967.4,-2844.1,-13903.,-1711.0,-1399.7,-5291.8,-2964.5,-5765.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
620.0000000000,6610.2,1377.7,1576.6,1337.3,1888.8,870.62,2244.8,337.78,1225.5,235.61,506.39,643.10,0.0000,-3920.7,-6911.1,-343.80,-2966.3,-2840.7,-13902.,-1710.1,-1395.6,-5290.5,-2963.7,-5763.9,1180.6,527.70,404.23,379.38,735.45,253.43,908.42,262.51,401.31,119.79,172.16,207.37,0.0000,-1.2800,-1.3318,-0.19112,-1.1788,-0.90977,-4.6546,-3.7557,-0.38225,-3.3678,-0.43042,-4.6691
621.0000000000,6580.8,1370.6,1587.5,1344.3,1885.9,903.61,2242.9,339.01,1239.8,237.75,506.21,645.69,0.0000,-3960.6,-6926.8,-346.87,-2965.8,-2866.2,-13902.,-1711.3,-1417.2,-5301.3,-2965.7,-5771.2,13687.,6118.0,4686.5,4398.5,8526.6,2938.2,10532.,3043.5,4652.7,1388.8,1995.9,2404.2,0.0000,-14.868,-15.447,-2.2158,-13.684,-10.578,-53.967,-43.542,-4.4317,-39.044,-4.9897,-54.130
622.0000000000,6575.7,1367.8,1585.1,1341.9,1874.3,909.43,2246.9,338.85,1246.1,237.44,511.94,649.18,0.0000,-3979.3,-6944.9,-349.89,-2965.3,-2874.5,-13901.,-1711.8,-1429.4,-5304.4,-2966.3,-5773.7,10785.,4820.5,3692.6,3465.7,6718.3,2315.1,8298.4,2398.0,3666.0,1094.3,1572.6,1894.3,0.0000,-11.741,-12.182,-1.7459,-10.793,-8.3521,-42.524,-34.308,-3.4918,-30.764,-3.9319,-42.650
623.0000000000,6652.6,1359.5,1574.4,1337.2,1874.9,893.93,2248.7,340.73,1234.1,239.07,511.95,647.92,0.0000,-3947.2,-6938.4,-348.15,-2964.6,-2852.3,-13900.,-1710.8,-1412.3,-5293.7,-2963.7,-5766.3,1004.2,448.87,343.84,322.71,625.59,215.57,772.72,223.30,341.37,101.89,146.44,176.39,0.0000,-1.0924,-1.1342,-0.16257,-1.0042,-0.77626,-3.9597,-3.1946,-0.32515,-2.8646,-0.36604,-3.9713
624.0000000000,6740.7,1353.3,1567.5,1335.9,1883.5,888.15,2256.7,341.46,1230.7,239.67,511.76,646.06,0.0000,-3935.6,-6928.4,-346.14,-2963.5,-2846.4,-13899.,-1709.8,-1404.5,-5290.2,-2962.5,-5763.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
625.0000000000,6822.8,1349.1,1565.3,1346.0,1912.4,900.67,2262.5,341.27,1237.1,241.39,509.53,643.18,0.0000,-3973.5,-6942.2,-348.60,-2962.4,-2870.3,-13899.,-1710.2,-1424.8,-5300.4,-2964.2,-5770.1,8031.0,3589.7,2749.8,2580.8,5003.0,1724.0,6179.6,1785.8,2730.0,814.87,1171.1,1410.7,0.0000,-8.7420,-9.0698,-1.3002,-8.0332,-6.2094,-31.664,-25.547,-2.6003,-22.908,-2.9261,-31.755
626.0000000000,6834.9,1338.8,1553.1,1343.5,1908.7,890.52,2262.3,340.28,1238.5,241.96,505.07,639.20,0.0000,-3943.4,-6934.7,-347.04,-2961.1,-2849.7,-13897.,-1709.5,-1410.0,-5291.6,-2961.7,-5763.8,200.90,89.797,68.787,64.559,125.15,43.126,154.58,44.671,68.291,20.384,29.295,35.288,0.0000,-0.21845,-0.22681,-0.32523E-01,-0.20079,-0.15502,-0.79200,-0.63903,-0.65046E-01,-0.57302,-0.73170E-01,-0.79428
627.0000000000,6851.0,1348.6,1561.5,1347.9,1934.2,903.23,2266.0,341.15,1246.0,241.10,504.40,641.46,0.0000,-3978.9,-6947.7,-349.37,-2960.2,-2872.3,-13897.,-1720.0,-1428.6,-5302.5,-2963.0,-5772.2,82542.,36895.,28262.,26525.,51420.,17719.,63513.,18354.,28058.,8375.1,12036.,14499.,0.0000,-89.905,-93.237,-13.363,-82.574,-63.814,-325.38,-262.57,-26.725,-235.43,-30.058,-326.32
628.0000000000,6883.5,1355.0,1560.2,1354.2,1803.4,896.52,2269.1,342.87,1249.0,239.50,508.15,640.07,0.0000,-3995.2,-6962.9,-351.77,-2959.5,-2879.5,-13896.,-1717.8,-1439.0,-5305.9,-2963.4,-5775.2,7216.7,3225.7,2471.0,2319.1,4495.7,1549.2,5553.0,1604.7,2453.2,732.24,1052.4,1267.6,0.0000,-7.8751,-8.1583,-1.1683,-7.2252,-5.5884,-28.446,-22.956,-2.3366,-20.584,-2.6277,-28.529
629.0000000000,6907.0,1346.1,1559.4,1353.4,1805.3,895.25,2291.6,343.13,1254.2,238.09,510.05,639.62,0.0000,-4008.4,-6977.3,-353.73,-2958.8,-2884.8,-13896.,-1720.4,-1446.8,-5307.6,-2963.4,-5777.1,40440.,18076.,13847.,12996.,25193.,8681.3,31118.,8992.2,13747.,4103.3,5897.2,7103.4,0.0000,-44.213,-45.759,-6.5469,-40.516,-31.360,-159.41,-128.64,-13.094,-115.35,-14.723,-159.86
630.0000000000,6951.6,1344.1,1575.8,1357.1,1807.3,899.68,2319.7,342.65,1256.0,237.66,513.43,643.14,0.0000,-4020.1,-6990.3,-355.29,-2958.0,-2889.9,-13895.,-1720.2,-1453.4,-5308.4,-2963.3,-5778.2,24020.,10737.,8224.5,7719.0,14964.,5156.4,18483.,5341.1,8165.2,2437.2,3502.7,4219.2,0.0000,-26.310,-27.207,-3.8887,-24.082,-18.656,-94.682,-76.412,-7.7773,-68.513,-8.7435,-94.957
631.0000000000,6967.5,1347.1,1550.5,1360.5,1838.8,890.70,2330.6,342.38,1240.8,236.27,516.65,644.76,0.0000,-3984.4,-6978.3,-352.44,-2957.1,-2866.9,-13894.,-1716.6,-1432.3,-5296.5,-2960.7,-5769.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
632.0000000000,6974.2,1347.1,1512.9,1358.1,1852.2,890.71,2331.7,343.39,1227.4,236.18,518.42,644.30,0.0000,-3970.2,-6964.4,-349.65,-2955.8,-2860.2,-13894.,-1713.9,-1422.2,-5292.2,-2959.5,-5766.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
633.0000000000,6983.7,1342.8,1513.3,1366.4,1874.2,897.41,2340.3,344.22,1228.6,239.25,523.12,646.51,0.0000,-3959.8,-6951.1,-347.46,-2954.6,-2855.7,-13894.,-1712.0,-1415.3,-5290.2,-2958.6,-5763.6,835.03,373.24,285.91,268.34,520.19,179.25,642.53,185.67,283.85,84.726,121.77,146.67,0.0000,-0.91209,-0.94481,-0.13518,-0.83541,-0.64558,-3.2928,-2.6568,-0.27037,-2.3820,-0.30390,-3.3020
634.0000000000,7003.8,1340.0,1527.8,1376.8,1882.2,909.93,2336.1,343.05,1231.9,240.66,528.37,648.39,0.0000,-3997.5,-6963.2,-349.91,-2953.8,-2879.9,-13895.,-1710.9,-1435.6,-5300.5,-2960.5,-5769.8,2087.6,933.13,714.81,670.87,1300.5,448.15,1606.4,464.20,709.65,211.82,304.43,366.70,0.0000,-2.2841,-2.3629,-0.33797,-2.0908,-1.6178,-8.2325,-6.6423,-0.67594,-5.9553,-0.75975,-8.2559
635.0000000000,7028.6,1348.0,1531.1,1384.0,1878.7,918.15,2332.6,344.93,1236.7,237.99,532.98,651.50,0.0000,-4014.0,-6977.8,-352.49,-2953.4,-2887.2,-13895.,-1734.1,-1446.2,-5308.3,-2961.3,-5777.6,0.18009E+06,80497.,61663.,57873.,0.11219E+06,38660.,0.13857E+06,40044.,61218.,18273.,26261.,31633.,0.0000,-197.38,-203.97,-29.155,-180.51,-139.80,-710.17,-573.12,-58.310,-513.75,-65.537,-712.24
636.0000000000,7022.5,1350.8,1534.4,1385.8,1882.6,919.70,2336.7,346.04,1252.3,235.40,533.89,655.98,0.0000,-4026.8,-6991.1,-354.58,-2952.9,-2892.6,-13895.,-1731.6,-1453.8,-5312.1,-2961.6,-5781.9,31677.,14159.,10846.,10180.,19734.,6800.1,24375.,7043.7,10768.,3214.1,4619.3,5564.2,0.0000,-34.780,-35.909,-5.1283,-31.776,-24.625,-124.93,-100.82,-10.257,-90.371,-11.526,-125.31
637.0000000000,7037.7,1397.7,1556.3,1378.7,1905.1,953.77,2395.1,356.66,1240.0,243.74,553.19,668.85,0.0000,-3993.5,-6980.8,-352.13,-2953.0,-2871.3,-13897.,-1725.0,-1433.1,-5301.3,-2960.7,-5774.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
638.0000000000,7043.2,1398.3,1560.2,1376.4,1937.5,920.34,2359.6,353.06,1227.6,243.15,557.79,663.92,0.0000,-3980.5,-6968.4,-349.64,-2952.5,-2864.7,-13898.,-1719.9,-1423.4,-5298.1,-2961.2,-5770.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
639.0000000000,7064.5,1407.7,1544.4,1381.5,1944.2,911.78,2347.5,354.89,1230.4,241.34,566.30,671.34,0.0000,-3970.4,-6954.9,-347.67,-2951.9,-2859.9,-13898.,-1716.2,-1416.4,-5295.6,-2962.1,-5767.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
640.0000000000,7127.9,1416.6,1553.6,1372.8,1935.0,906.72,2369.3,355.57,1222.9,242.48,580.29,664.38,0.0000,-3961.4,-6944.2,-346.19,-2950.8,-2855.9,-13898.,-1713.5,-1411.0,-5293.6,-2963.8,-5764.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
641.0000000000,7148.7,1433.7,1545.6,1370.5,1959.8,902.12,2359.6,364.69,1234.7,240.96,598.69,667.04,0.0000,-3952.7,-6935.3,-345.04,-2949.5,-2852.0,-13898.,-1711.7,-1406.4,-5292.0,-2966.0,-5763.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
642.0000000000,7193.0,1432.5,1527.8,1370.4,1959.3,906.14,2353.0,363.25,1233.2,241.45,590.65,668.49,0.0000,-3945.5,-6926.3,-344.11,-2948.1,-2848.2,-13898.,-1710.3,-1402.3,-5290.5,-2966.9,-5761.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
643.0000000000,7383.2,1434.5,1518.0,1369.6,1948.0,899.59,2370.3,361.68,1241.3,240.62,581.55,663.39,0.0000,-3939.0,-6917.4,-343.32,-2946.8,-2844.3,-13897.,-1709.4,-1398.7,-5288.9,-2966.3,-5760.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
644.0000000000,7412.0,1424.4,1519.6,1371.2,1937.7,897.96,2373.5,358.74,1258.5,238.97,577.67,657.66,0.0000,-3932.0,-6909.5,-342.63,-2945.2,-2840.6,-13898.,-1708.7,-1395.4,-5287.4,-2965.4,-5759.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
645.0000000000,7420.4,1425.8,1521.7,1372.9,1952.6,897.36,2388.2,359.75,1260.2,239.58,571.47,653.42,0.0000,-3925.7,-6901.9,-342.01,-2943.5,-2837.1,-13898.,-1708.2,-1392.6,-5286.2,-2964.5,-5758.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
646.0000000000,7418.5,1422.9,1533.8,1380.3,1965.7,897.09,2392.3,358.17,1263.1,239.69,565.10,651.64,0.0000,-3919.8,-6895.2,-341.45,-2942.1,-2833.7,-13898.,-1707.8,-1390.0,-5285.2,-2963.4,-5758.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
647.0000000000,7404.8,1418.9,1540.0,1385.1,1959.8,904.38,2400.5,358.40,1257.5,240.16,562.89,651.20,0.0000,-3914.5,-6889.5,-340.93,-2940.7,-2830.4,-13898.,-1707.5,-1387.5,-5284.3,-2962.2,-5757.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
648.0000000000,7392.3,1404.1,1546.9,1384.7,1964.2,911.08,2402.4,356.18,1252.7,242.52,559.92,647.72,0.0000,-3909.0,-6884.4,-340.42,-2939.5,-2827.2,-13898.,-1707.3,-1385.2,-5283.5,-2960.7,-5757.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
649.0000000000,7393.5,1399.5,1554.6,1388.9,1974.3,928.88,2400.4,358.38,1257.2,242.80,564.98,646.59,0.0000,-3949.8,-6902.8,-344.05,-2938.7,-2852.2,-13899.,-1717.2,-1407.8,-5296.5,-2961.8,-5767.9,74652.,33368.,25561.,23990.,46505.,16025.,57442.,16599.,25376.,7574.6,10886.,13113.,0.0000,-80.989,-84.000,-12.085,-74.515,-57.140,-294.27,-237.66,-24.171,-213.00,-27.106,-295.32
650.0000000000,7392.8,1393.7,1535.0,1384.1,1971.5,916.03,2403.1,358.25,1241.0,241.15,570.02,644.47,0.0000,-3921.7,-6899.6,-343.34,-2938.0,-2832.2,-13898.,-1714.6,-1395.8,-5289.1,-2959.4,-5763.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
651.0000000000,7394.8,1382.3,1533.0,1374.9,1957.3,907.73,2396.2,358.08,1230.1,242.10,574.16,648.14,0.0000,-3911.5,-6892.3,-342.13,-2937.5,-2827.2,-13898.,-1712.4,-1390.6,-5286.7,-2959.0,-5761.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
652.0000000000,7351.9,1376.7,1532.9,1377.5,1945.8,905.10,2394.2,357.29,1246.2,242.35,572.95,649.80,0.0000,-3903.8,-6885.3,-341.04,-2936.9,-2823.7,-13897.,-1710.7,-1387.1,-5285.3,-2958.4,-5760.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
653.0000000000,7366.5,1373.2,1531.9,1385.4,1940.7,897.83,2402.2,357.13,1253.3,242.39,575.83,646.74,0.0000,-3896.9,-6879.5,-340.12,-2936.3,-2820.6,-13896.,-1709.5,-1384.4,-5284.2,-2957.7,-5760.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
654.0000000000,7380.4,1373.1,1535.1,1394.5,1964.0,898.64,2391.8,355.94,1263.7,242.47,570.95,646.03,0.0000,-3890.8,-6873.9,-339.34,-2935.4,-2817.6,-13896.,-1708.6,-1382.3,-5283.1,-2956.8,-5759.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
655.0000000000,7376.3,1377.7,1540.8,1396.9,1968.2,908.23,2394.7,355.58,1264.2,245.64,574.05,641.86,0.0000,-3885.3,-6868.5,-338.66,-2934.7,-2815.2,-13895.,-1707.9,-1380.2,-5282.3,-2956.0,-5758.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
656.0000000000,7381.2,1379.4,1540.5,1397.6,1979.5,908.15,2409.6,355.38,1266.0,244.46,575.61,637.04,0.0000,-3880.4,-6863.9,-338.05,-2934.4,-2812.7,-13895.,-1707.5,-1378.3,-5282.0,-2955.4,-5757.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
657.0000000000,7373.0,1369.9,1533.5,1399.2,1973.0,906.49,2398.8,353.91,1276.5,245.76,570.79,634.76,0.0000,-3875.4,-6860.4,-337.50,-2933.9,-2810.1,-13895.,-1707.1,-1376.5,-5281.7,-2954.3,-5756.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
658.0000000000,7370.8,1363.2,1524.2,1398.1,1982.1,907.79,2385.7,353.51,1277.7,245.31,566.98,634.97,0.0000,-3870.7,-6856.6,-336.98,-2933.3,-2807.6,-13894.,-1706.8,-1374.9,-5281.2,-2953.4,-5756.1,5.5359,2.4744,1.8955,1.7790,3.4486,1.1884,4.2597,1.2309,1.8818,0.56170,0.80726,0.97239,0.0000,-0.59527E-02,-0.61986E-02,-0.89621E-03,-0.55042E-02,-0.41901E-02,-0.21817E-01,-0.17616E-01,-0.17924E-02,-0.15791E-01,-0.20059E-02,-0.21877E-01
659.0000000000,7374.2,1378.4,1524.7,1406.4,1988.8,941.39,2380.3,354.65,1284.4,245.63,563.02,638.57,0.0000,-3912.4,-6877.3,-340.60,-2933.0,-2833.3,-13894.,-1707.1,-1397.3,-5292.2,-2955.1,-5763.4,3088.3,1380.4,1057.4,992.43,1923.9,662.95,2376.3,686.70,1049.8,313.35,450.34,542.46,0.0000,-3.3271,-3.4594,-0.49996,-3.0744,-2.3436,-12.170,-9.8266,-0.99992,-8.8092,-1.1189,-12.203
660.0000000000,7220.0,1344.3,1526.2,1406.7,1988.1,937.86,2377.6,355.84,1283.6,245.16,562.26,639.30,0.0000,-3932.3,-6899.6,-344.02,-2933.0,-2842.0,-13894.,-1708.8,-1410.9,-5295.7,-2955.6,-5766.1,14104.,6304.4,4829.3,4532.5,8786.4,3027.8,10853.,3136.2,4794.5,1431.1,2056.8,2477.5,0.0000,-15.228,-15.813,-2.2834,-14.056,-10.727,-55.582,-44.877,-4.5668,-40.232,-5.1093,-55.727
661.0000000000,7195.7,1337.3,1518.8,1403.3,1990.8,945.67,2351.6,357.37,1286.3,243.57,563.84,642.28,0.0000,-3948.3,-6919.8,-346.72,-2933.5,-2848.9,-13894.,-1713.9,-1421.3,-5297.9,-2955.8,-5768.6,42401.,18952.,14518.,13626.,26414.,9102.1,32626.,9428.1,14413.,4302.2,6183.0,7447.8,0.0000,-45.878,-47.583,-6.8643,-42.291,-32.307,-167.09,-134.91,-13.729,-120.94,-15.358,-167.51
662.0000000000,7196.7,1324.2,1496.7,1402.8,1982.3,929.07,2351.2,358.07,1277.0,244.97,568.15,643.74,0.0000,-3915.6,-6914.0,-344.69,-2933.5,-2826.7,-13893.,-1711.9,-1404.3,-5287.1,-2953.4,-5761.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
663.0000000000,7198.1,1317.2,1505.3,1401.7,1987.6,926.21,2343.7,356.38,1286.7,245.75,572.16,644.32,0.0000,-3903.6,-6904.2,-342.47,-2933.3,-2821.0,-13892.,-1710.3,-1396.9,-5283.6,-2952.5,-5758.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
664.0000000000,7193.7,1309.3,1499.8,1402.6,1971.1,918.65,2336.3,353.27,1288.2,245.01,570.46,647.45,0.0000,-3894.8,-6894.2,-340.68,-2932.8,-2817.2,-13891.,-1709.0,-1391.9,-5281.7,-2951.8,-5757.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
665.0000000000,7194.0,1316.7,1490.1,1404.6,1971.2,913.20,2340.1,350.66,1288.8,243.68,567.10,646.03,0.0000,-3887.3,-6885.1,-339.29,-2932.0,-2813.9,-13891.,-1708.1,-1388.0,-5280.4,-2951.3,-5755.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
666.0000000000,7195.3,1334.4,1486.7,1416.4,1976.8,903.76,2347.9,348.91,1287.5,243.13,565.98,642.65,0.0000,-3880.4,-6877.2,-338.20,-2931.0,-2810.8,-13890.,-1707.4,-1384.6,-5279.3,-2950.6,-5754.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
667.0000000000,7304.7,1349.2,1491.5,1407.6,1984.4,902.47,2358.8,346.72,1284.8,243.42,567.11,643.85,0.0000,-3874.2,-6870.3,-337.31,-2930.1,-2807.8,-13889.,-1706.9,-1381.6,-5278.3,-2949.6,-5753.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
668.0000000000,7318.5,1361.3,1501.2,1405.9,1994.3,901.62,2363.0,343.79,1291.0,242.82,564.50,647.75,0.0000,-3868.3,-6864.1,-336.56,-2929.2,-2804.9,-13889.,-1706.5,-1379.1,-5277.5,-2948.8,-5752.8,0.65058,0.29080,0.22276,0.20907,0.40528,0.13966,0.50060,0.14466,0.22115,0.66011E-01,0.94870E-01,0.11428,0.0000,-0.69899E-03,-0.72740E-03,-0.10532E-03,-0.64635E-03,-0.49039E-03,-0.25630E-02,-0.20693E-02,-0.21065E-03,-0.18553E-02,-0.23526E-03,-0.25682E-02
669.0000000000,7317.8,1350.4,1499.9,1401.8,1986.1,901.63,2358.6,347.38,1291.4,242.58,566.36,650.17,0.0000,-3862.7,-6858.4,-335.91,-2928.2,-2802.2,-13888.,-1706.2,-1376.8,-5276.7,-2947.9,-5752.0,0.65058,0.29080,0.22276,0.20907,0.40528,0.13966,0.50060,0.14466,0.22115,0.66011E-01,0.94870E-01,0.11428,0.0000,-0.69835E-03,-0.72690E-03,-0.10532E-03,-0.64609E-03,-0.48971E-03,-0.25629E-02,-0.20692E-02,-0.21065E-03,-0.18552E-02,-0.23520E-03,-0.25679E-02
670.0000000000,7318.0,1344.3,1498.0,1402.1,1982.2,901.88,2362.3,345.89,1292.4,243.29,569.14,649.67,0.0000,-3857.3,-6853.1,-335.33,-2927.4,-2799.6,-13887.,-1706.0,-1374.7,-5276.1,-2947.1,-5751.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
671.0000000000,7315.6,1344.5,1486.8,1403.1,1964.1,897.63,2361.0,343.58,1279.6,243.33,569.91,647.60,0.0000,-3852.0,-6848.1,-334.81,-2926.5,-2797.1,-13887.,-1705.8,-1372.6,-5275.5,-2946.4,-5750.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
672.0000000000,7307.3,1347.5,1477.9,1407.3,1961.0,900.23,2355.9,343.83,1282.7,242.25,572.45,647.30,0.0000,-3847.1,-6843.6,-334.32,-2925.7,-2794.6,-13886.,-1705.7,-1370.7,-5275.0,-2945.7,-5749.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
673.0000000000,7294.3,1343.2,1469.2,1409.6,1957.6,901.38,2353.4,346.36,1266.9,241.15,572.35,645.02,0.0000,-3842.1,-6839.3,-333.86,-2924.8,-2792.1,-13885.,-1705.6,-1369.0,-5274.3,-2945.2,-5749.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
674.0000000000,7295.2,1347.0,1479.2,1418.5,1941.5,916.23,2353.2,347.85,1277.2,240.29,569.45,644.14,0.0000,-3883.3,-6858.7,-337.53,-2924.1,-2817.7,-13885.,-1739.3,-1391.2,-5292.2,-2947.2,-5765.7,0.25088E+06,0.11214E+06,85903.,80623.,0.15629E+06,53857.,0.19305E+06,55786.,85283.,25456.,36585.,44068.,0.0000,-268.80,-279.68,-40.616,-249.11,-188.43,-987.99,-797.95,-81.232,-715.35,-90.610,-989.72
675.0000000000,7325.1,1344.4,1489.9,1425.4,1931.8,933.01,2375.8,351.67,1275.2,242.73,568.97,654.69,0.0000,-3903.0,-6879.6,-340.99,-2923.8,-2826.9,-13886.,-1749.6,-1404.9,-5302.5,-2947.9,-5777.4,0.13896E+06,62113.,47580.,44656.,86567.,29830.,0.10693E+06,30899.,47237.,14100.,20264.,24409.,0.0000,-149.20,-155.07,-22.497,-138.15,-104.65,-547.37,-442.09,-44.993,-396.25,-50.183,-548.35
676.0000000000,7339.4,1439.9,1546.6,1431.1,1977.1,1025.5,2488.0,363.98,1264.8,261.14,605.12,688.18,0.0000,-3923.9,-6901.9,-343.83,-2925.1,-2838.4,-13890.,-1738.7,-1415.4,-5306.5,-2950.8,-5781.0,4684.6,2093.9,1604.0,1505.4,2918.3,1005.6,3604.7,1041.7,1592.4,475.32,683.13,822.86,0.0000,-5.0576,-5.2393,-0.75840,-4.6699,-3.5548,-18.483,-14.913,-1.5168,-13.364,-1.6955,-18.509
677.0000000000,7338.8,1442.2,1553.4,1433.0,1969.1,992.19,2463.4,360.15,1272.3,268.37,617.05,688.32,0.0000,-3942.1,-6924.0,-346.10,-2926.4,-2845.6,-13894.,-1729.9,-1424.3,-5309.8,-2953.9,-5780.2,3162.2,1413.4,1082.7,1016.2,1969.9,678.81,2433.2,703.13,1074.9,320.85,461.12,555.44,0.0000,-3.4256,-3.5415,-0.51193,-3.1566,-2.4082,-12.484,-10.070,-1.0239,-9.0231,-1.1456,-12.503
678.0000000000,7342.6,1428.4,1509.0,1427.5,1980.5,939.06,2404.6,366.97,1282.8,259.20,619.70,697.11,0.0000,-3910.2,-6915.7,-343.78,-2927.1,-2822.2,-13894.,-1722.9,-1406.3,-5297.2,-2953.7,-5770.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
679.0000000000,7340.7,1404.7,1530.8,1430.0,1984.0,905.23,2398.3,366.50,1283.6,256.53,639.09,683.78,0.0000,-3898.3,-6905.8,-341.47,-2926.4,-2815.3,-13894.,-1717.8,-1398.4,-5291.9,-2955.5,-5765.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
680.0000000000,7374.7,1406.5,1517.0,1421.6,1999.6,893.92,2394.5,368.72,1294.4,253.18,645.24,679.79,0.0000,-3888.8,-6896.2,-339.69,-2924.9,-2810.8,-13894.,-1714.3,-1393.4,-5288.4,-2957.5,-5761.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
681.0000000000,7372.1,1399.3,1497.0,1425.7,2008.1,906.23,2398.8,373.15,1283.4,253.74,649.17,684.07,0.0000,-3881.7,-6887.5,-338.33,-2923.5,-2807.1,-13893.,-1711.8,-1389.5,-5285.6,-2958.9,-5759.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
682.0000000000,7360.1,1382.2,1499.9,1427.7,1987.7,922.03,2427.5,372.84,1279.4,253.75,631.61,678.97,0.0000,-3875.9,-6878.8,-337.28,-2922.0,-2803.6,-13893.,-1710.1,-1386.0,-5283.2,-2958.1,-5757.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
683.0000000000,7371.5,1367.9,1499.7,1429.1,1984.4,914.15,2461.4,366.96,1289.4,254.35,624.98,673.04,0.0000,-3870.1,-6871.1,-336.44,-2920.5,-2800.0,-13893.,-1708.9,-1383.0,-5281.3,-2957.0,-5755.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
684.0000000000,7382.0,1361.7,1489.2,1434.5,1997.0,913.32,2472.4,367.49,1278.5,256.59,609.22,675.67,0.0000,-3864.3,-6864.1,-335.72,-2919.2,-2796.7,-13893.,-1708.0,-1380.3,-5280.1,-2955.5,-5754.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
685.0000000000,7483.4,1358.5,1498.3,1424.8,1991.9,922.82,2470.6,363.46,1274.6,255.69,602.28,674.11,0.0000,-3859.0,-6857.3,-335.10,-2918.0,-2793.5,-13893.,-1707.4,-1377.8,-5279.0,-2953.9,-5753.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
686.0000000000,7579.8,1354.9,1511.2,1424.8,1996.0,923.63,2484.4,360.57,1279.4,256.06,594.15,674.77,0.0000,-3854.4,-6851.7,-334.54,-2917.0,-2790.5,-13893.,-1706.9,-1375.5,-5277.9,-2952.0,-5753.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
687.0000000000,7580.7,1335.9,1506.0,1423.9,2049.2,926.79,2485.1,360.45,1285.7,257.60,589.89,675.61,0.0000,-3849.4,-6846.7,-334.03,-2916.1,-2787.6,-13892.,-1706.5,-1373.4,-5277.2,-2950.5,-5752.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
688.0000000000,7579.7,1334.2,1508.3,1425.0,2049.0,925.47,2469.0,361.83,1284.9,257.94,591.41,676.75,0.0000,-3844.2,-6842.3,-333.56,-2915.3,-2785.0,-13892.,-1706.2,-1371.6,-5276.6,-2949.7,-5752.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
689.0000000000,7594.8,1325.7,1513.0,1429.2,2041.9,933.60,2447.7,356.35,1283.3,257.45,594.84,680.98,0.0000,-3839.2,-6838.5,-333.11,-2914.5,-2782.5,-13891.,-1706.0,-1369.8,-5276.0,-2949.5,-5752.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
690.0000000000,7659.0,1320.6,1516.4,1432.1,2034.2,937.90,2459.5,357.50,1292.3,258.48,595.80,688.02,0.0000,-3834.1,-6835.5,-332.67,-2913.8,-2780.1,-13890.,-1705.9,-1368.2,-5276.0,-2949.5,-5751.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
691.0000000000,7729.1,1325.0,1523.7,1439.9,2026.1,938.40,2460.3,359.00,1297.8,257.60,596.33,690.40,0.0000,-3829.2,-6832.2,-332.25,-2913.2,-2777.7,-13889.,-1705.7,-1367.1,-5275.7,-2949.3,-5751.6,35.355,15.803,12.105,11.361,22.024,7.5895,27.204,7.8613,12.018,3.5873,5.1555,6.2101,0.0000,-0.37723E-01,-0.39270E-01,-0.57236E-02,-0.35019E-01,-0.26282E-01,-0.13926,-0.11253,-0.11447E-01,-0.10086,-0.12751E-01,-0.13962
692.0000000000,7725.1,1344.2,1526.5,1452.3,2033.4,964.31,2473.4,357.81,1309.5,259.51,594.43,690.11,0.0000,-3871.3,-6852.4,-335.93,-2912.9,-2803.6,-13890.,-1708.7,-1389.7,-5287.5,-2951.5,-5760.0,22585.,10095.,7733.1,7257.7,14069.,4848.2,17378.,5021.9,7677.3,2291.6,3293.4,3967.1,0.0000,-24.138,-25.099,-3.6563,-22.399,-16.834,-88.960,-71.885,-7.3126,-64.427,-8.1446,-89.175
693.0000000000,7718.4,1336.3,1526.3,1459.9,2047.2,957.43,2488.8,357.82,1302.2,262.97,591.41,686.09,0.0000,-3845.4,-6850.7,-335.28,-2913.0,-2784.4,-13889.,-1707.8,-1379.2,-5280.1,-2948.7,-5754.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
694.0000000000,7731.2,1340.3,1519.6,1458.6,2052.3,963.71,2479.8,355.86,1322.7,262.70,595.41,678.26,0.0000,-3837.6,-6845.1,-334.13,-2913.1,-2780.0,-13889.,-1707.1,-1374.8,-5277.7,-2947.1,-5752.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
695.0000000000,7747.6,1328.6,1516.2,1455.3,2040.3,960.34,2476.9,353.18,1335.6,262.30,591.93,674.37,0.0000,-3832.3,-6839.8,-333.11,-2913.1,-2777.2,-13888.,-1706.5,-1371.7,-5276.5,-2945.6,-5751.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
696.0000000000,7754.4,1337.8,1508.9,1455.5,2021.0,970.87,2467.3,353.17,1338.0,261.14,587.49,676.93,0.0000,-3827.5,-6835.7,-332.27,-2912.7,-2774.5,-13887.,-1706.1,-1369.2,-5275.3,-2944.3,-5750.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
697.0000000000,7774.6,1332.8,1487.1,1454.6,2028.4,969.47,2465.0,353.81,1332.0,258.56,581.44,677.60,0.0000,-3823.0,-6831.8,-331.56,-2912.6,-2772.5,-13887.,-1705.8,-1367.2,-5274.0,-2943.0,-5749.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
698.0000000000,7724.0,1327.6,1481.5,1460.2,2053.0,964.19,2469.0,351.51,1331.3,260.41,590.31,684.04,0.0000,-3818.3,-6827.9,-330.95,-2912.4,-2770.6,-13887.,-1705.5,-1365.4,-5273.2,-2942.5,-5749.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
699.0000000000,7606.8,1332.1,1457.3,1465.3,2053.6,949.45,2473.9,349.50,1337.6,258.67,592.41,683.13,0.0000,-3813.8,-6823.4,-330.42,-2912.1,-2768.6,-13886.,-1705.3,-1363.8,-5272.6,-2942.2,-5748.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
700.0000000000,7620.4,1339.8,1454.4,1469.3,2050.5,948.91,2472.0,350.30,1322.6,258.55,592.62,681.17,0.0000,-3809.3,-6819.4,-329.94,-2911.3,-2766.2,-13886.,-1705.2,-1362.3,-5272.0,-2941.7,-5747.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
701.0000000000,7661.9,1363.3,1453.8,1469.6,2062.4,952.84,2488.2,349.99,1316.9,257.02,588.43,682.33,0.0000,-3805.0,-6815.8,-329.50,-2910.4,-2764.0,-13885.,-1705.0,-1361.1,-5271.4,-2940.9,-5747.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
702.0000000000,7756.8,1330.5,1462.2,1474.1,2061.0,961.68,2491.8,354.83,1331.2,257.58,595.04,687.03,0.0000,-3800.9,-6812.5,-329.07,-2909.7,-2761.9,-13885.,-1704.9,-1360.0,-5271.0,-2940.2,-5747.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
703.0000000000,7764.5,1299.7,1458.6,1484.1,2034.0,965.63,2479.4,352.89,1329.0,255.48,593.09,689.64,0.0000,-3796.8,-6809.5,-328.67,-2909.1,-2759.9,-13884.,-1704.8,-1358.9,-5270.4,-2939.4,-5746.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
704.0000000000,7781.5,1279.3,1459.5,1487.4,2039.9,982.25,2468.0,355.13,1326.7,255.97,582.92,689.16,0.0000,-3792.9,-6806.7,-328.28,-2908.5,-2757.9,-13884.,-1704.7,-1357.9,-5269.9,-2938.7,-5746.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
705.0000000000,7794.4,1262.1,1463.7,1482.2,2048.2,981.02,2456.9,352.92,1334.2,257.37,588.13,686.31,0.0000,-3788.8,-6804.5,-327.91,-2908.0,-2756.1,-13883.,-1704.6,-1357.0,-5269.5,-2938.1,-5745.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
706.0000000000,7819.0,1263.3,1454.8,1481.0,2053.2,969.84,2462.5,350.66,1333.8,256.44,590.22,685.88,0.0000,-3785.0,-6803.2,-327.54,-2907.5,-2754.2,-13881.,-1704.5,-1356.0,-5269.2,-2937.6,-5745.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
707.0000000000,7821.8,1272.2,1439.2,1487.9,2034.5,968.38,2446.2,349.31,1334.9,256.01,586.79,686.77,0.0000,-3781.3,-6800.6,-327.18,-2907.0,-2752.4,-13880.,-1704.5,-1355.0,-5268.9,-2937.1,-5744.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
708.0000000000,7824.2,1275.5,1431.0,1488.9,2021.7,958.71,2454.0,346.69,1346.6,255.51,584.43,688.69,0.0000,-3777.7,-6798.2,-326.82,-2906.3,-2750.5,-13879.,-1704.4,-1354.1,-5268.6,-2936.5,-5744.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
709.0000000000,7809.3,1268.0,1436.0,1487.8,2034.0,955.40,2435.0,341.97,1360.3,254.29,591.35,688.06,0.0000,-3774.1,-6795.8,-326.48,-2905.7,-2748.6,-13878.,-1704.3,-1353.1,-5268.2,-2935.9,-5743.7,306.72,137.10,105.02,98.565,191.07,65.843,236.01,68.201,104.26,31.121,44.727,53.876,0.0000,-0.32400,-0.33785,-0.49655E-01,-0.30243,-0.22426,-1.2070,-0.97509,-0.99310E-01,-0.87435,-0.11017,-1.2078
710.0000000000,7804.2,1260.2,1436.0,1488.0,2033.9,958.53,2413.9,340.88,1363.8,253.84,586.70,686.13,0.0000,-3770.7,-6793.6,-326.14,-2905.0,-2746.8,-13877.,-1704.4,-1352.1,-5267.9,-2935.0,-5743.3,1316.3,588.35,450.69,422.99,819.99,282.56,1012.8,292.68,447.44,133.56,191.94,231.21,0.0000,-1.3895,-1.4491,-0.21309,-1.2975,-0.96134,-5.1797,-4.1843,-0.42619,-3.7521,-0.47271,-5.1825
711.0000000000,7804.3,1257.3,1438.4,1491.4,2037.8,960.13,2406.4,342.04,1365.8,252.38,585.78,684.44,0.0000,-3767.3,-6791.3,-325.81,-2904.3,-2744.9,-13876.,-1704.3,-1351.2,-5267.5,-2934.2,-5742.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
712.0000000000,7809.5,1262.9,1438.7,1496.2,2036.7,964.25,2429.7,341.17,1373.8,250.30,587.96,684.34,0.0000,-3764.1,-6788.9,-325.49,-2903.6,-2743.1,-13876.,-1704.2,-1350.4,-5267.0,-2933.4,-5742.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
713.0000000000,7898.1,1253.0,1435.7,1501.7,2040.0,967.29,2433.2,339.01,1370.9,250.01,587.11,685.73,0.0000,-3760.8,-6786.5,-325.17,-2902.9,-2741.3,-13875.,-1704.1,-1349.5,-5266.5,-2932.8,-5741.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
714.0000000000,7922.9,1241.6,1429.2,1503.1,2028.2,967.90,2428.8,338.31,1371.8,251.37,582.56,684.96,0.0000,-3757.6,-6784.4,-324.86,-2902.2,-2739.5,-13874.,-1704.0,-1348.4,-5266.2,-2932.1,-5741.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
715.0000000000,8043.8,1243.9,1422.6,1505.5,2017.4,969.21,2427.1,339.13,1375.1,252.08,583.82,684.49,0.0000,-3754.2,-6782.4,-324.55,-2901.5,-2737.8,-13873.,-1703.9,-1347.5,-5265.8,-2931.6,-5740.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
716.0000000000,8147.3,1237.2,1415.2,1502.7,2018.2,967.73,2407.1,340.12,1376.9,250.74,585.16,685.12,0.0000,-3750.8,-6780.5,-324.25,-2900.8,-2736.0,-13872.,-1703.8,-1346.6,-5265.3,-2931.0,-5740.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
717.0000000000,8111.0,1226.9,1403.8,1499.1,2018.8,972.01,2403.6,341.22,1380.7,249.87,585.45,686.03,0.0000,-3747.5,-6778.5,-323.95,-2899.8,-2734.2,-13871.,-1703.7,-1345.7,-5264.7,-2930.4,-5739.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
718.0000000000,8124.9,1217.9,1412.9,1510.0,2011.4,986.29,2411.0,342.21,1387.3,249.01,583.68,686.03,0.0000,-3789.6,-6799.9,-327.74,-2899.0,-2760.5,-13872.,-1704.0,-1367.2,-5275.6,-2932.5,-5747.4,2556.9,1142.9,875.48,821.67,1592.8,548.88,1967.4,568.54,869.17,259.44,372.85,449.12,0.0000,-2.6926,-2.8063,-0.41394,-2.5192,-1.8590,-10.057,-8.1238,-0.82788,-7.2865,-0.91701,-10.056
719.0000000000,8287.8,1205.4,1406.3,1502.1,2002.7,983.24,2418.1,344.69,1375.9,248.95,584.95,684.98,0.0000,-3764.7,-6799.7,-327.24,-2898.0,-2741.7,-13871.,-1703.9,-1358.0,-5267.2,-2930.5,-5741.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
720.0000000000,8381.1,1200.6,1400.9,1500.6,1995.6,981.01,2428.9,343.17,1377.2,250.09,586.55,684.51,0.0000,-3757.5,-6795.8,-326.22,-2896.9,-2737.7,-13870.,-1703.7,-1354.3,-5264.7,-2929.6,-5740.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
721.0000000000,8383.7,1197.7,1399.7,1511.6,2003.8,978.83,2418.2,343.80,1377.1,250.23,586.64,682.02,0.0000,-3752.4,-6791.4,-325.33,-2895.8,-2735.1,-13869.,-1703.6,-1352.1,-5263.7,-2928.9,-5739.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
722.0000000000,8464.4,1200.5,1393.4,1520.7,2000.7,991.94,2419.2,341.99,1383.9,250.15,581.91,681.97,0.0000,-3793.2,-6810.3,-328.68,-2895.1,-2760.9,-13870.,-1703.8,-1373.2,-5274.6,-2931.0,-5746.5,2431.3,1086.7,832.47,781.30,1514.6,521.92,1870.8,540.61,826.47,246.69,354.54,427.06,0.0000,-2.5610,-2.6677,-0.39360,-2.3954,-1.7650,-9.5608,-7.7229,-0.78720,-6.9277,-0.87145,-9.5567
723.0000000000,8536.2,1201.9,1392.1,1526.4,1999.3,995.23,2425.8,341.86,1378.7,250.71,578.38,681.19,0.0000,-3812.8,-6831.4,-331.96,-2894.4,-2769.9,-13869.,-1704.1,-1386.6,-5277.7,-2931.6,-5749.0,3068.3,1371.5,1050.6,986.01,1911.4,658.67,2361.0,682.26,1043.0,311.33,447.43,538.95,0.0000,-3.2388,-3.3700,-0.49673,-3.0262,-2.2324,-12.065,-9.7458,-0.99346,-8.7426,-1.0997,-12.059
724.0000000000,8589.5,1196.1,1383.9,1519.4,1999.2,972.54,2431.8,340.65,1373.2,248.40,579.91,679.76,0.0000,-3783.0,-6827.6,-330.51,-2893.3,-2748.4,-13868.,-1703.9,-1372.8,-5267.4,-2929.2,-5742.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
725.0000000000,8547.2,1189.9,1362.0,1516.6,2001.3,962.69,2433.0,341.04,1376.4,245.01,575.58,681.19,0.0000,-3773.3,-6820.1,-328.73,-2892.1,-2743.2,-13866.,-1703.6,-1366.8,-5264.2,-2927.9,-5739.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
726.0000000000,8569.4,1183.6,1352.9,1517.4,1998.6,961.86,2428.3,341.35,1382.2,245.13,577.05,684.68,0.0000,-3766.7,-6812.7,-327.28,-2890.9,-2740.0,-13865.,-1703.4,-1363.1,-5262.8,-2926.9,-5738.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
727.0000000000,8574.8,1187.7,1359.0,1531.0,1997.3,976.57,2420.2,336.90,1402.4,244.83,578.69,687.40,0.0000,-3806.4,-6829.2,-330.24,-2890.0,-2765.3,-13865.,-1716.3,-1383.6,-5276.1,-2928.6,-5749.2,96879.,43303.,33171.,31132.,60351.,20797.,74545.,21542.,32932.,9829.8,14127.,17017.,0.0000,-102.26,-106.38,-15.684,-95.486,-70.302,-380.84,-307.68,-31.367,-276.01,-34.701,-380.57
728.0000000000,8585.8,1177.7,1382.1,1544.6,1994.7,986.92,2422.6,335.76,1420.5,245.71,578.17,691.21,0.0000,-3825.1,-6848.0,-333.23,-2889.4,-2773.9,-13865.,-1713.6,-1396.1,-5280.4,-2929.0,-5753.2,4327.5,1934.3,1481.7,1390.7,2695.9,928.98,3329.9,962.26,1471.1,439.09,631.06,760.14,0.0000,-4.5770,-4.7564,-0.70059,-4.2695,-3.1470,-17.011,-13.744,-1.4012,-12.329,-1.5500,-16.998
729.0000000000,8578.4,1173.5,1385.7,1547.4,1984.7,972.72,2423.1,333.86,1432.5,248.22,581.34,694.92,0.0000,-3794.3,-6842.0,-331.56,-2888.6,-2752.3,-13863.,-1710.6,-1381.0,-5269.9,-2926.5,-5746.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
730.0000000000,8578.0,1176.3,1390.2,1542.3,1964.6,989.22,2415.1,331.96,1449.5,248.95,588.90,697.19,0.0000,-3829.7,-6856.1,-333.72,-2888.1,-2774.9,-13863.,-1709.1,-1398.5,-5277.9,-2927.9,-5751.1,5575.9,2492.3,1909.2,1791.8,3473.5,1197.0,4290.4,1239.8,1895.4,565.75,813.09,979.41,0.0000,-5.9049,-6.1328,-0.90268,-5.5021,-4.0551,-21.915,-17.707,-1.8054,-15.885,-1.9965,-21.897
731.0000000000,8578.0,1177.3,1390.6,1547.0,1956.0,995.77,2406.4,332.96,1450.3,249.16,590.34,695.94,0.0000,-3846.2,-6872.1,-336.03,-2887.8,-2782.4,-13862.,-1709.8,-1409.1,-5280.0,-2928.1,-5752.7,18385.,8217.6,6294.9,5908.0,11453.,3946.6,14146.,4088.0,6249.5,1865.4,2680.9,3229.3,0.0000,-19.506,-20.240,-2.9763,-18.157,-13.395,-72.255,-58.382,-5.9526,-52.375,-6.5821,-72.194
732.0000000000,8593.4,1169.0,1393.1,1551.5,1961.4,997.56,2408.8,332.59,1434.8,250.94,589.54,694.74,0.0000,-3859.7,-6887.1,-337.96,-2887.4,-2788.1,-13862.,-1711.8,-1417.2,-5281.2,-2928.2,-5753.9,29372.,13129.,10057.,9438.8,18297.,6305.2,22601.,6531.1,9984.4,2980.2,4283.1,5159.2,0.0000,-31.224,-32.371,-4.7550,-29.029,-21.435,-115.43,-93.271,-9.5101,-83.675,-10.515,-115.33
733.0000000000,8594.5,1160.8,1394.9,1560.1,1965.9,999.97,2414.1,333.32,1434.2,251.18,589.45,696.34,0.0000,-3872.1,-6900.6,-339.55,-2887.0,-2793.4,-13861.,-1713.9,-1424.2,-5282.2,-2928.1,-5755.1,33244.,14859.,11383.,10683.,20710.,7136.4,25580.,7392.0,11301.,3373.1,4847.7,5839.4,0.0000,-35.407,-36.679,-5.3819,-32.880,-24.299,-130.64,-105.57,-10.764,-94.706,-11.899,-130.53
734.0000000000,8544.5,1156.2,1387.6,1554.8,1965.0,989.38,2422.7,331.76,1426.2,251.73,587.64,697.28,0.0000,-3837.3,-6889.3,-336.77,-2886.4,-2770.4,-13859.,-1710.9,-1404.6,-5270.8,-2925.4,-5747.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
735.0000000000,8548.8,1161.9,1377.1,1555.8,1964.7,984.43,2432.9,329.97,1423.1,251.89,589.06,701.23,0.0000,-3824.2,-6875.1,-334.04,-2885.5,-2764.2,-13858.,-1708.5,-1395.1,-5266.6,-2924.2,-5743.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
736.0000000000,8599.6,1134.1,1371.4,1556.1,1967.9,985.59,2432.3,332.27,1427.2,251.01,585.97,707.48,0.0000,-3814.6,-6862.1,-331.91,-2884.4,-2759.9,-13858.,-1706.7,-1388.6,-5264.3,-2923.2,-5741.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
737.0000000000,8644.0,1127.2,1372.3,1560.8,1967.3,995.65,2432.7,335.94,1433.3,251.98,586.69,708.02,0.0000,-3806.6,-6850.4,-330.30,-2883.5,-2756.7,-13857.,-1705.5,-1383.4,-5262.9,-2922.6,-5739.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
738.0000000000,8641.5,1127.9,1370.0,1566.4,1955.3,995.59,2430.2,336.90,1438.0,251.30,586.41,710.69,0.0000,-3799.6,-6839.9,-329.07,-2882.5,-2753.5,-13857.,-1704.5,-1378.9,-5262.0,-2922.1,-5738.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
739.0000000000,8584.9,1131.7,1375.8,1568.0,1953.5,1014.0,2437.4,335.54,1451.7,252.06,586.51,707.35,0.0000,-3838.8,-6854.4,-332.19,-2881.7,-2778.5,-13857.,-1704.2,-1399.4,-5273.0,-2924.2,-5745.1,2192.4,979.97,750.68,704.54,1365.8,470.64,1687.0,487.50,745.27,222.45,319.71,385.10,0.0000,-2.3298,-2.4147,-0.35493,-2.1643,-1.5953,-8.6184,-6.9628,-0.70987,-6.2463,-0.78415,-8.6097
740.0000000000,8455.5,1124.6,1378.7,1570.5,1950.8,1023.8,2433.1,336.30,1455.1,250.35,585.77,705.15,0.0000,-3856.6,-6871.4,-335.27,-2881.1,-2786.5,-13857.,-1710.0,-1411.1,-5277.1,-2924.7,-5748.6,46754.,20898.,16009.,15025.,29126.,10037.,35976.,10396.,15893.,4743.9,6817.8,8212.4,0.0000,-49.770,-51.534,-7.5690,-46.197,-34.083,-183.78,-148.49,-15.138,-133.20,-16.720,-183.60
741.0000000000,8486.1,1120.9,1378.4,1575.2,1953.5,1030.9,2428.4,335.80,1458.1,249.92,586.44,698.84,0.0000,-3870.7,-6887.1,-337.67,-2880.8,-2792.2,-13857.,-1708.7,-1419.7,-5278.8,-2925.1,-5750.0,4786.4,2139.4,1638.9,1538.1,2981.7,1027.5,3683.0,1064.3,1627.0,485.65,697.97,840.74,0.0000,-5.1039,-5.2805,-0.77487,-4.7329,-3.4948,-18.813,-15.201,-1.5497,-13.636,-1.7113,-18.795
742.0000000000,8521.6,1114.3,1366.1,1571.4,1952.9,1019.1,2428.1,335.68,1455.9,246.88,591.21,704.57,0.0000,-3837.0,-6877.4,-335.42,-2880.1,-2769.2,-13855.,-1707.0,-1401.2,-5267.6,-2922.6,-5742.1,171.91,76.841,58.863,55.245,107.09,36.904,132.28,38.226,58.438,17.443,25.069,30.197,0.0000,-0.18320,-0.18964,-0.27831E-01,-0.16984,-0.12522,-0.67567,-0.54597,-0.55662E-01,-0.48977,-0.61447E-01,-0.67503
743.0000000000,8533.6,1112.4,1371.3,1574.9,1961.1,1020.6,2438.8,335.78,1456.2,245.87,589.69,703.48,0.0000,-3824.3,-6864.5,-333.02,-2879.2,-2763.0,-13854.,-1705.6,-1392.5,-5263.6,-2921.4,-5739.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
744.0000000000,8525.7,1111.0,1362.0,1572.0,1961.5,1013.9,2450.2,334.82,1462.0,245.65,591.41,700.42,0.0000,-3814.9,-6852.4,-331.08,-2878.1,-2758.8,-13853.,-1704.5,-1386.6,-5261.5,-2920.3,-5737.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
745.0000000000,8525.9,1111.2,1359.9,1579.0,1961.1,1005.9,2445.7,336.71,1454.3,245.11,591.81,696.20,0.0000,-3806.8,-6841.5,-329.57,-2876.8,-2755.2,-13852.,-1703.7,-1381.8,-5260.1,-2919.6,-5735.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
746.0000000000,8525.2,1114.4,1353.2,1570.4,1948.4,1006.1,2455.9,335.85,1452.0,245.30,594.63,698.43,0.0000,-3799.5,-6832.0,-328.38,-2875.5,-2751.8,-13851.,-1703.2,-1377.8,-5259.1,-2919.0,-5734.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
747.0000000000,8567.9,1115.8,1347.5,1581.9,1951.8,1002.6,2468.4,336.33,1448.2,247.39,597.18,699.25,0.0000,-3792.6,-6823.8,-327.41,-2874.3,-2748.7,-13850.,-1702.7,-1374.2,-5258.3,-2918.6,-5733.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
748.0000000000,8680.9,1122.4,1333.2,1600.4,1954.6,1000.1,2478.3,335.35,1451.7,248.46,600.02,699.60,0.0000,-3786.3,-6815.8,-326.60,-2873.2,-2745.9,-13848.,-1702.4,-1371.1,-5257.6,-2918.3,-5732.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
749.0000000000,8673.4,1125.3,1327.2,1601.4,1954.9,993.56,2494.2,332.77,1446.7,246.84,603.54,700.04,0.0000,-3780.7,-6808.4,-325.88,-2872.1,-2743.2,-13847.,-1702.2,-1368.2,-5256.9,-2917.9,-5731.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
750.0000000000,8725.7,1122.8,1315.6,1596.4,1952.0,990.06,2495.5,333.43,1436.3,247.98,605.98,701.31,0.0000,-3775.2,-6802.3,-325.24,-2870.9,-2740.3,-13846.,-1702.0,-1365.6,-5256.2,-2917.5,-5730.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
751.0000000000,8816.0,1117.3,1307.3,1584.7,1961.3,997.78,2509.1,335.88,1435.6,247.97,607.24,702.18,0.0000,-3769.8,-6796.8,-324.65,-2869.8,-2737.5,-13845.,-1701.8,-1363.1,-5255.7,-2917.2,-5730.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
752.0000000000,8818.6,1119.5,1308.8,1597.2,1959.6,1018.2,2502.1,334.12,1442.9,248.75,605.39,703.24,0.0000,-3810.3,-6814.7,-328.19,-2869.0,-2763.0,-13845.,-1705.9,-1384.4,-5267.6,-2919.4,-5738.5,31008.,13860.,10617.,9964.5,19317.,6656.4,23860.,6894.9,10541.,3146.2,4521.7,5446.6,0.0000,-32.809,-34.006,-5.0199,-30.538,-22.331,-121.82,-98.444,-10.040,-88.323,-11.055,-121.65
753.0000000000,8830.1,1121.1,1317.0,1597.8,1954.5,1029.8,2474.5,333.89,1440.7,249.93,605.55,702.06,0.0000,-3829.5,-6834.7,-331.54,-2868.5,-2771.5,-13843.,-1709.6,-1397.4,-5272.2,-2920.1,-5742.4,35745.,15977.,12239.,11487.,22267.,7673.2,27504.,7948.1,12151.,3626.8,5212.4,6278.6,0.0000,-37.890,-39.232,-5.7867,-35.240,-25.796,-140.43,-113.48,-11.573,-101.81,-12.741,-140.22
754.0000000000,8830.9,1117.8,1320.7,1596.7,1957.6,1026.7,2476.9,333.25,1439.5,249.92,605.52,703.45,0.0000,-3844.7,-6853.2,-334.18,-2867.9,-2777.7,-13842.,-1707.8,-1407.2,-5273.7,-2920.3,-5743.9,2259.8,1010.1,773.76,726.20,1407.8,485.11,1738.9,502.49,768.18,229.29,329.53,396.94,0.0000,-2.4000,-2.4827,-0.36584,-2.2299,-1.6337,-8.8779,-7.1743,-0.73169,-6.4367,-0.80539,-8.8642
755.0000000000,8830.7,1116.9,1312.2,1581.1,1960.5,1013.5,2490.0,333.76,1445.0,249.38,604.85,699.98,0.0000,-3812.3,-6846.0,-332.13,-2867.2,-2755.1,-13840.,-1706.0,-1390.2,-5262.5,-2917.9,-5736.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
756.0000000000,8830.5,1117.1,1312.8,1577.8,1963.2,1018.6,2502.7,334.34,1440.1,248.58,605.27,695.80,0.0000,-3800.6,-6835.3,-329.87,-2866.1,-2749.1,-13838.,-1704.6,-1382.4,-5258.8,-2916.7,-5732.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
757.0000000000,8825.1,1104.7,1308.2,1570.3,1968.8,1016.1,2513.5,333.89,1436.1,248.77,606.83,695.11,0.0000,-3792.0,-6825.2,-328.04,-2865.0,-2745.0,-13837.,-1703.5,-1377.0,-5256.9,-2915.7,-5731.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
758.0000000000,8815.5,1093.6,1309.4,1569.6,1974.3,1008.8,2520.8,331.87,1428.1,248.19,607.76,697.60,0.0000,-3784.7,-6816.2,-326.61,-2863.9,-2741.6,-13836.,-1702.7,-1372.7,-5255.6,-2914.9,-5729.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
759.0000000000,8824.5,1086.5,1292.3,1573.4,1972.9,999.67,2531.5,332.04,1432.7,248.87,609.00,700.67,0.0000,-3778.1,-6808.1,-325.47,-2862.8,-2738.6,-13835.,-1702.2,-1369.1,-5254.6,-2914.2,-5728.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
760.0000000000,8863.0,1078.4,1287.3,1579.0,1979.7,993.21,2550.1,331.88,1428.0,250.31,612.67,696.38,0.0000,-3772.0,-6800.9,-324.55,-2861.7,-2736.0,-13834.,-1701.8,-1365.9,-5253.8,-2913.6,-5727.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
761.0000000000,8955.0,1072.3,1275.2,1599.3,2007.2,1008.1,2559.6,332.14,1434.4,249.69,613.68,693.64,0.0000,-3812.3,-6817.6,-327.86,-2861.1,-2761.5,-13835.,-1705.3,-1386.7,-5265.4,-2915.7,-5735.6,28252.,12628.,9673.3,9078.8,17600.,6064.7,21739.,6282.0,9603.6,2866.6,4119.7,4962.4,0.0000,-29.894,-30.955,-4.5737,-27.815,-20.271,-110.98,-89.671,-9.1474,-80.459,-10.051,-110.77
762.0000000000,8947.7,1067.5,1278.6,1606.5,2018.8,1011.1,2561.5,333.25,1427.6,248.05,615.08,694.65,0.0000,-3831.1,-6837.1,-331.06,-2860.5,-2769.9,-13834.,-1709.4,-1399.0,-5269.9,-2916.2,-5739.5,39097.,17476.,13387.,12564.,24356.,8392.8,30084.,8693.5,13290.,3967.0,5701.2,6867.5,0.0000,-41.445,-42.873,-6.3294,-38.531,-28.111,-153.59,-124.10,-12.659,-111.35,-13.907,-153.29
763.0000000000,8934.7,1049.4,1270.6,1602.8,1973.1,996.47,2561.9,334.28,1416.9,247.61,615.87,698.02,0.0000,-3799.9,-6831.5,-329.53,-2859.7,-2748.0,-13833.,-1707.2,-1383.4,-5260.0,-2913.8,-5732.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
764.0000000000,8969.2,1041.6,1268.3,1595.1,1825.0,989.58,2568.4,335.12,1415.3,247.62,616.37,699.96,0.0000,-3789.0,-6821.9,-327.65,-2858.7,-2742.3,-13833.,-1705.3,-1376.2,-5256.8,-2912.6,-5729.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
765.0000000000,9073.4,1045.2,1258.2,1594.9,1828.7,1006.7,2579.3,336.10,1429.1,248.65,616.05,699.62,0.0000,-3826.9,-6836.0,-330.20,-2858.0,-2766.6,-13833.,-1704.2,-1395.6,-5266.5,-2914.2,-5735.9,1928.2,861.89,660.23,619.65,1201.2,413.93,1483.7,428.76,655.47,195.65,281.18,338.70,0.0000,-2.0440,-2.1143,-0.31217,-1.8996,-1.3841,-7.5745,-6.1199,-0.62433,-5.4913,-0.68534,-7.5591
766.0000000000,9072.4,1031.6,1253.0,1566.1,1830.9,995.51,2591.6,336.53,1431.4,247.27,614.71,700.38,0.0000,-3798.1,-6829.1,-328.76,-2857.2,-2746.3,-13832.,-1703.1,-1382.0,-5257.3,-2912.0,-5729.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
767.0000000000,9068.6,1035.9,1246.3,1560.1,1832.7,995.90,2599.2,335.94,1428.0,247.49,614.77,704.40,0.0000,-3787.9,-6819.7,-327.05,-2856.3,-2741.2,-13831.,-1702.3,-1375.4,-5254.3,-2911.0,-5726.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
768.0000000000,9074.2,1031.6,1248.2,1562.4,1829.1,997.88,2606.6,336.23,1424.3,248.31,617.05,707.74,0.0000,-3780.3,-6810.6,-325.63,-2855.2,-2737.8,-13830.,-1701.7,-1370.7,-5252.8,-2910.2,-5725.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
769.0000000000,9087.8,1027.5,1251.3,1561.1,1832.3,993.03,2613.6,336.24,1427.4,245.74,614.64,712.43,0.0000,-3773.5,-6802.5,-324.50,-2853.9,-2734.7,-13830.,-1701.2,-1366.9,-5251.8,-2909.4,-5724.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
770.0000000000,9098.6,1020.9,1233.3,1557.3,1840.1,992.50,2602.0,336.24,1426.0,246.33,610.94,712.25,0.0000,-3767.4,-6795.2,-323.58,-2852.7,-2731.9,-13829.,-1700.9,-1363.6,-5251.1,-2908.9,-5723.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
771.0000000000,9078.5,1017.6,1176.4,1553.4,1846.2,982.76,2596.0,335.53,1427.2,246.16,608.91,713.98,0.0000,-3761.6,-6788.5,-322.82,-2851.5,-2729.2,-13828.,-1700.6,-1360.6,-5250.6,-2908.4,-5722.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
772.0000000000,9082.6,1018.4,1174.6,1564.7,1848.7,976.02,2589.2,337.44,1433.4,247.12,608.88,716.26,0.0000,-3756.1,-6782.7,-322.16,-2850.4,-2726.5,-13828.,-1700.4,-1358.0,-5250.2,-2907.9,-5721.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
773.0000000000,9085.3,1017.1,1173.4,1565.1,1852.8,970.14,2599.0,337.70,1433.0,246.62,608.36,711.99,0.0000,-3750.9,-6777.1,-321.58,-2849.4,-2723.9,-13827.,-1700.2,-1355.6,-5249.8,-2907.5,-5720.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
774.0000000000,9092.7,1018.1,1164.1,1566.2,1854.9,961.14,2604.3,338.41,1436.4,247.01,611.87,712.82,0.0000,-3745.9,-6772.0,-321.05,-2848.3,-2721.3,-13826.,-1700.0,-1353.4,-5249.4,-2907.1,-5720.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
775.0000000000,9093.9,1018.6,1157.4,1566.7,1853.6,965.67,2594.4,339.19,1443.4,247.98,614.42,709.14,0.0000,-3741.0,-6767.2,-320.55,-2847.3,-2718.9,-13825.,-1699.9,-1351.3,-5249.1,-2906.9,-5719.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
776.0000000000,9113.3,1018.1,1157.5,1569.6,1851.3,959.94,2587.9,338.79,1449.0,248.65,615.19,709.10,0.0000,-3736.3,-6762.6,-320.08,-2846.2,-2716.5,-13824.,-1699.8,-1349.4,-5248.7,-2906.5,-5719.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
777.0000000000,9211.7,1009.1,1149.6,1565.7,1838.1,950.17,2587.0,337.56,1458.3,247.76,613.02,708.72,0.0000,-3731.7,-6758.4,-319.63,-2845.2,-2714.2,-13823.,-1699.7,-1347.6,-5248.1,-2906.2,-5718.8,626.18,279.89,214.40,201.22,390.08,134.42,481.82,139.24,212.86,63.535,91.312,109.99,0.0000,-0.65686,-0.68157,-0.10137,-0.61365,-0.44216,-2.4591,-1.9865,-0.20275,-1.7829,-0.22190,-2.4530
778.0000000000,9223.6,1008.7,1146.7,1560.4,1832.0,964.96,2600.3,337.20,1462.9,247.31,612.59,708.58,0.0000,-3772.6,-6778.0,-323.29,-2844.6,-2740.0,-13823.,-1700.1,-1368.6,-5259.1,-2908.5,-5726.4,3137.3,1402.3,1074.2,1008.2,1954.4,673.47,2414.0,697.59,1066.5,318.32,457.49,551.07,0.0000,-3.2964,-3.4163,-0.50789,-3.0785,-2.2214,-12.320,-9.9523,-1.0158,-8.9322,-1.1117,-12.289
779.0000000000,9224.9,999.81,1139.2,1548.5,1831.6,958.89,2603.5,338.18,1453.1,246.92,607.51,708.74,0.0000,-3746.6,-6775.7,-322.68,-2843.8,-2720.8,-13822.,-1699.9,-1358.4,-5250.8,-2906.8,-5720.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
780.0000000000,9225.7,996.46,1128.0,1548.5,1831.3,958.18,2616.3,338.79,1444.4,246.21,609.05,708.41,0.0000,-3738.4,-6769.9,-321.56,-2842.8,-2716.3,-13821.,-1699.7,-1354.0,-5248.4,-2906.1,-5719.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
781.0000000000,9249.2,974.48,1126.1,1558.4,1839.8,959.96,2618.9,337.04,1449.2,246.05,611.63,709.36,0.0000,-3732.6,-6763.8,-320.58,-2841.8,-2713.4,-13820.,-1699.5,-1351.2,-5247.4,-2905.5,-5718.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
782.0000000000,9269.0,960.46,1123.9,1561.0,1855.5,962.29,2618.5,337.35,1450.8,244.98,612.66,706.75,0.0000,-3727.4,-6758.3,-319.77,-2840.8,-2710.8,-13819.,-1699.4,-1349.0,-5246.7,-2905.0,-5717.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
783.0000000000,9271.9,965.21,1119.6,1561.3,1855.8,958.90,2606.9,337.63,1457.5,244.20,613.20,706.94,0.0000,-3722.6,-6753.2,-319.09,-2839.8,-2708.3,-13819.,-1699.2,-1347.1,-5246.2,-2904.6,-5717.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
784.0000000000,9233.1,969.81,1220.1,1563.1,1851.6,963.39,2593.8,337.48,1460.7,244.11,616.08,705.15,0.0000,-3718.2,-6748.6,-318.51,-2838.8,-2705.9,-13818.,-1699.1,-1345.3,-5245.7,-2904.2,-5716.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
785.0000000000,9082.7,968.97,1223.2,1562.6,1843.4,960.88,2593.9,336.18,1476.8,244.29,617.93,702.27,0.0000,-3713.9,-6744.5,-318.00,-2837.8,-2703.6,-13818.,-1699.0,-1343.7,-5245.3,-2903.7,-5716.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
786.0000000000,9102.5,971.61,1220.7,1555.1,1812.3,950.54,2598.6,333.74,1482.0,245.86,619.10,701.39,0.0000,-3709.8,-6740.7,-317.53,-2836.9,-2701.4,-13817.,-1698.9,-1342.3,-5245.0,-2903.2,-5716.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
787.0000000000,9117.0,978.20,1225.6,1550.2,1815.9,957.40,2592.2,335.01,1478.0,247.18,614.74,696.76,0.0000,-3705.9,-6736.8,-317.09,-2836.0,-2699.2,-13816.,-1698.7,-1340.9,-5244.7,-2902.6,-5715.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
788.0000000000,9104.5,988.01,1226.7,1560.3,1808.7,963.49,2612.0,337.60,1491.9,247.40,614.54,699.56,0.0000,-3702.1,-6733.3,-316.68,-2835.2,-2697.1,-13816.,-1698.6,-1339.6,-5244.4,-2901.8,-5715.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
789.0000000000,9103.5,992.11,1233.4,1567.2,1803.4,981.85,2589.8,334.93,1504.6,246.87,615.01,699.21,0.0000,-3743.5,-6753.3,-320.35,-2834.7,-2723.0,-13815.,-1700.2,-1360.5,-5255.9,-2903.7,-5723.5,11661.,5212.1,3992.6,3747.2,7264.2,2503.2,8972.6,2592.9,3963.9,1183.2,1700.4,2048.2,0.0000,-12.184,-12.648,-1.8878,-11.414,-8.1692,-45.780,-36.971,-3.7755,-33.190,-4.1191,-45.638
790.0000000000,9117.4,997.13,1232.5,1572.2,1799.4,985.87,2590.1,333.56,1505.8,247.99,612.43,699.68,0.0000,-3763.6,-6775.4,-323.85,-2834.5,-2732.0,-13815.,-1700.2,-1374.1,-5259.5,-2904.1,-5726.3,3319.0,1483.5,1136.4,1066.6,2067.6,712.48,2553.9,738.00,1128.2,336.76,483.99,582.99,0.0000,-3.4750,-3.6016,-0.53732,-3.2524,-2.3307,-13.030,-10.522,-1.0746,-9.4467,-1.1722,-12.989
791.0000000000,9149.8,1005.2,1234.1,1573.1,1801.7,989.34,2591.0,330.05,1508.2,249.98,615.31,702.62,0.0000,-3780.0,-6795.5,-326.65,-2834.2,-2738.8,-13814.,-1700.0,-1384.6,-5260.8,-2904.1,-5727.4,1378.1,615.96,471.84,442.84,858.46,295.82,1060.4,306.42,468.44,139.82,200.95,242.06,0.0000,-1.4459,-1.4963,-0.22309,-1.3517,-0.96968,-5.4100,-4.3687,-0.44619,-3.9222,-0.48664,-5.3927
792.0000000000,9179.6,1008.9,1228.9,1551.8,1795.3,972.37,2586.1,325.52,1501.0,249.24,612.29,700.57,0.0000,-3749.2,-6789.8,-324.75,-2833.7,-2716.7,-13813.,-1699.5,-1369.3,-5249.8,-2901.3,-5719.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
793.0000000000,9181.8,1007.1,1214.2,1548.0,1793.6,959.57,2564.9,321.78,1500.0,249.73,612.72,702.04,0.0000,-3738.9,-6780.7,-322.64,-2832.9,-2711.1,-13811.,-1699.1,-1362.5,-5246.5,-2899.8,-5717.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
794.0000000000,9146.0,1002.9,1218.3,1550.9,1799.1,964.08,2564.8,320.66,1512.6,250.94,613.20,704.63,0.0000,-3776.9,-6795.1,-325.02,-2832.4,-2735.6,-13811.,-1704.5,-1381.6,-5257.8,-2901.4,-5725.4,42843.,19150.,14669.,13768.,26689.,9197.0,32966.,9526.5,14564.,4347.1,6247.5,7525.4,0.0000,-44.976,-46.533,-6.9359,-42.006,-30.097,-168.18,-135.81,-13.872,-121.93,-15.118,-167.62
795.0000000000,9137.3,992.29,1204.8,1546.1,1803.9,956.59,2566.6,323.46,1496.8,249.79,614.15,698.67,0.0000,-3748.7,-6788.8,-323.51,-2831.7,-2715.6,-13809.,-1702.9,-1368.7,-5249.7,-2899.1,-5720.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
796.0000000000,9123.6,994.71,1205.5,1548.1,1803.9,949.17,2560.4,323.62,1490.2,249.32,611.14,698.36,0.0000,-3738.9,-6779.7,-321.77,-2830.9,-2710.7,-13808.,-1701.5,-1362.4,-5247.1,-2898.0,-5718.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
797.0000000000,8961.5,1001.0,1214.2,1548.6,1811.2,952.62,2546.9,324.48,1494.1,250.31,608.50,698.47,0.0000,-3777.0,-6794.2,-324.43,-2830.6,-2735.5,-13807.,-1702.3,-1381.8,-5257.6,-2899.8,-5725.2,13996.,6255.8,4792.1,4497.5,8718.7,3004.4,10769.,3112.0,4757.5,1420.1,2040.9,2458.4,0.0000,-14.693,-15.201,-2.2658,-13.719,-9.8218,-54.930,-44.359,-4.5315,-39.829,-4.9347,-54.743
798.0000000000,8949.3,1005.4,1219.6,1553.5,1810.4,960.43,2541.6,325.07,1490.5,251.23,610.60,696.50,0.0000,-3794.3,-6811.4,-327.20,-2830.4,-2743.8,-13806.,-1701.5,-1393.3,-5260.4,-2900.4,-5727.3,3201.2,1430.9,1096.1,1028.7,1994.2,687.19,2463.2,711.80,1088.2,324.81,466.81,562.29,0.0000,-3.3668,-3.4787,-0.51824,-3.1410,-2.2514,-12.563,-10.146,-1.0365,-9.1097,-1.1285,-12.520
799.0000000000,8958.8,1007.8,1218.2,1560.5,1807.9,964.33,2532.5,325.70,1494.7,250.68,610.99,693.48,0.0000,-3808.2,-6827.3,-329.47,-2830.3,-2750.0,-13804.,-1701.3,-1402.0,-5261.5,-2900.8,-5728.0,5619.7,2511.9,1924.2,1805.9,3500.8,1206.4,4324.1,1249.6,1910.3,570.20,819.48,987.10,0.0000,-5.9214,-6.1122,-0.90977,-5.5186,-3.9599,-22.054,-17.810,-1.8195,-15.992,-1.9807,-21.978
800.0000000000,8981.6,989.26,1207.0,1556.7,1812.4,945.35,2545.2,324.90,1479.0,247.43,611.42,693.92,0.0000,-3775.0,-6817.8,-327.19,-2829.8,-2727.5,-13802.,-1700.3,-1384.2,-5250.2,-2898.3,-5720.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
801.0000000000,8991.8,989.61,1203.6,1551.1,1816.7,936.48,2548.9,322.37,1473.9,248.03,609.93,696.29,0.0000,-3762.6,-6805.2,-324.80,-2829.1,-2721.4,-13800.,-1699.5,-1375.8,-5246.5,-2897.2,-5717.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
802.0000000000,9024.8,988.37,1200.7,1553.9,1823.4,932.86,2553.9,320.09,1465.8,248.14,610.95,698.94,0.0000,-3753.5,-6793.3,-322.89,-2828.2,-2717.4,-13798.,-1698.8,-1370.1,-5244.7,-2896.3,-5715.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
803.0000000000,9035.3,984.94,1211.2,1559.4,1818.2,933.55,2561.0,318.38,1449.1,247.36,614.97,698.59,0.0000,-3745.6,-6782.7,-321.43,-2827.3,-2714.1,-13796.,-1698.4,-1365.5,-5243.6,-2895.5,-5714.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
804.0000000000,9018.4,986.61,1215.1,1556.4,1815.1,929.20,2561.6,318.03,1438.2,247.98,615.57,698.38,0.0000,-3738.6,-6773.3,-320.29,-2826.4,-2711.0,-13795.,-1698.0,-1361.6,-5242.8,-2894.9,-5713.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
805.0000000000,9103.8,978.96,1213.7,1557.9,1818.6,926.10,2563.4,317.76,1435.0,248.52,617.49,696.86,0.0000,-3732.1,-6764.8,-319.38,-2825.6,-2708.2,-13793.,-1697.7,-1358.1,-5242.2,-2894.2,-5712.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
806.0000000000,9126.3,978.24,1211.8,1555.2,1821.9,917.55,2579.7,318.41,1434.1,249.59,619.36,698.90,0.0000,-3726.0,-6757.2,-318.62,-2824.8,-2705.5,-13792.,-1697.5,-1355.0,-5241.6,-2893.6,-5711.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
807.0000000000,9130.6,983.49,1215.9,1552.5,1810.8,923.30,2596.0,316.94,1455.3,250.80,623.86,702.10,0.0000,-3765.6,-6773.5,-322.02,-2824.3,-2731.0,-13791.,-1698.6,-1375.4,-5252.9,-2895.8,-5719.6,9187.7,4106.7,3145.9,2952.5,5723.6,1972.3,7069.7,2043.0,3123.2,932.24,1339.8,1613.8,0.0000,-9.6342,-9.9734,-1.4874,-8.9986,-6.4224,-36.052,-29.105,-2.9748,-26.140,-3.2313,-35.914
808.0000000000,9187.2,977.85,1213.5,1549.4,1825.5,913.40,2604.7,315.41,1448.8,250.57,623.33,700.96,0.0000,-3738.5,-6768.9,-321.22,-2823.8,-2711.6,-13789.,-1698.3,-1363.8,-5245.0,-2893.8,-5714.0,931.22,416.24,318.85,299.25,580.11,199.90,716.54,207.06,316.55,94.486,135.79,163.57,0.0000,-0.97591,-1.0107,-0.15076,-0.91155,-0.64989,-3.6540,-2.9498,-0.30151,-2.6493,-0.32742,-3.6399
809.0000000000,9189.9,989.33,1219.8,1544.0,1831.6,932.64,2614.8,312.73,1452.0,252.13,624.67,699.86,0.0000,-3774.9,-6784.6,-324.04,-2823.6,-2735.0,-13788.,-1704.4,-1382.0,-5255.6,-2895.6,-5721.7,48045.,21475.,16451.,15440.,29930.,10314.,36969.,10683.,16332.,4874.9,7006.1,8439.3,0.0000,-50.436,-52.164,-7.7781,-47.086,-33.618,-188.52,-152.20,-15.556,-136.69,-16.891,-187.79
810.0000000000,9172.0,994.37,1223.0,1541.8,1829.9,948.12,2612.0,313.29,1457.5,254.33,625.47,702.81,0.0000,-3792.1,-6802.0,-326.82,-2823.5,-2743.0,-13787.,-1725.9,-1393.1,-5263.7,-2896.2,-5730.5,0.17442E+06,77964.,59722.,56051.,0.10866E+06,37443.,0.13421E+06,38784.,59292.,17698.,25435.,30638.,0.0000,-183.45,-189.48,-28.237,-171.11,-122.31,-684.41,-552.64,-56.475,-496.24,-61.315,-681.74
811.0000000000,9169.7,995.45,1225.1,1538.0,1814.1,954.48,2638.6,314.34,1455.0,257.43,625.53,710.21,0.0000,-3806.1,-6818.3,-329.07,-2823.3,-2749.1,-13787.,-1732.0,-1401.7,-5269.8,-2896.3,-5737.5,99743.,44583.,34152.,32053.,62136.,21412.,76749.,22179.,33906.,10120.,14545.,17520.,0.0000,-105.12,-108.44,-16.147,-97.942,-70.084,-391.47,-316.09,-32.295,-283.79,-35.058,-389.95
812.0000000000,9191.6,1051.6,1251.8,1530.6,1837.7,1010.7,2740.2,322.75,1453.9,265.50,644.96,733.94,0.0000,-3776.2,-6811.2,-326.84,-2824.0,-2730.0,-13788.,-1722.6,-1383.9,-5260.2,-2895.0,-5731.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
813.0000000000,9202.8,1052.4,1280.1,1517.6,1828.2,994.48,2747.9,322.48,1459.5,275.37,657.29,731.85,0.0000,-3767.4,-6802.8,-324.52,-2824.1,-2725.8,-13791.,-1715.3,-1375.5,-5258.0,-2895.6,-5726.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
814.0000000000,9200.5,1040.2,1269.6,1515.2,1822.9,962.33,2702.5,318.40,1453.2,271.21,649.08,722.54,0.0000,-3760.0,-6791.8,-322.68,-2824.1,-2721.5,-13792.,-1709.9,-1369.7,-5255.9,-2895.8,-5723.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
815.0000000000,9111.9,1039.9,1255.5,1528.6,1836.4,958.03,2664.3,323.33,1466.8,266.78,650.55,731.21,0.0000,-3798.5,-6804.0,-325.34,-2824.3,-2745.4,-13792.,-1706.9,-1389.2,-5265.1,-2898.2,-5728.4,6028.8,2694.8,2064.3,1937.4,3755.7,1294.2,4639.0,1340.5,2049.4,611.71,879.14,1059.0,0.0000,-6.3637,-6.5568,-0.97601,-5.9244,-4.2531,-23.703,-19.128,-1.9520,-17.165,-2.1219,-23.603
816.0000000000,9041.3,1037.1,1254.4,1529.8,1852.8,941.75,2671.9,325.21,1467.6,261.58,653.03,727.84,0.0000,-3770.2,-6796.1,-324.05,-2823.9,-2725.0,-13791.,-1704.0,-1375.7,-5255.0,-2897.2,-5720.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
817.0000000000,9015.1,1020.2,1272.3,1525.1,1866.6,933.87,2666.1,325.14,1473.0,261.25,662.00,720.78,0.0000,-3759.8,-6787.3,-322.51,-2823.0,-2719.4,-13790.,-1702.0,-1369.1,-5251.4,-2897.4,-5717.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
818.0000000000,8945.4,1022.7,1257.6,1515.8,1862.6,938.27,2661.3,325.29,1485.4,262.10,663.96,717.45,0.0000,-3751.5,-6778.1,-321.23,-2822.0,-2715.7,-13790.,-1700.5,-1364.5,-5249.5,-2898.0,-5714.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
819.0000000000,8848.9,1019.0,1243.5,1518.1,1829.3,937.75,2657.9,328.31,1480.5,258.31,666.89,722.60,0.0000,-3744.5,-6770.1,-320.22,-2821.2,-2712.3,-13789.,-1699.5,-1360.7,-5247.8,-2898.7,-5713.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
820.0000000000,8957.6,1006.0,1239.2,1514.1,1822.3,941.44,2661.5,330.44,1487.4,259.38,661.00,720.25,0.0000,-3738.8,-6762.0,-319.39,-2820.4,-2709.2,-13788.,-1698.7,-1357.4,-5246.3,-2898.2,-5712.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
821.0000000000,8947.2,997.51,1238.1,1517.4,1815.3,938.98,2671.0,332.62,1498.4,259.56,662.81,719.75,0.0000,-3733.1,-6754.8,-318.71,-2819.5,-2706.2,-13787.,-1698.2,-1354.4,-5245.1,-2897.4,-5711.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
822.0000000000,8937.7,991.34,1240.7,1517.2,1821.9,936.48,2689.5,331.97,1491.9,260.11,661.63,720.00,0.0000,-3727.8,-6748.5,-318.12,-2818.5,-2703.4,-13787.,-1697.7,-1351.7,-5244.0,-2896.8,-5710.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
823.0000000000,8952.8,997.06,1240.3,1518.0,1818.3,932.30,2696.9,331.94,1483.7,262.25,660.57,717.93,0.0000,-3722.7,-6742.8,-317.61,-2817.5,-2700.6,-13787.,-1697.4,-1349.2,-5243.1,-2896.3,-5709.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
824.0000000000,8977.2,992.20,1243.6,1513.5,1764.9,930.32,2715.0,332.93,1483.7,264.10,658.22,719.81,0.0000,-3718.0,-6737.1,-317.13,-2816.6,-2697.9,-13786.,-1697.2,-1346.9,-5242.6,-2895.5,-5708.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
825.0000000000,8993.4,989.66,1244.3,1505.7,1697.8,932.22,2711.8,329.19,1478.1,265.16,656.20,720.61,0.0000,-3713.5,-6731.9,-316.68,-2815.8,-2695.3,-13786.,-1697.0,-1344.8,-5242.0,-2894.5,-5708.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
826.0000000000,9014.1,986.49,1252.7,1509.9,1700.1,950.09,2711.9,328.86,1485.3,266.27,651.87,721.65,0.0000,-3754.7,-6751.0,-320.32,-2815.3,-2720.7,-13787.,-1698.0,-1365.4,-5253.2,-2895.9,-5716.4,8636.9,3860.5,2957.3,2775.5,5380.4,1854.1,6645.8,1920.5,2935.9,876.34,1259.5,1517.1,0.0000,-9.0378,-9.3575,-1.3982,-8.4565,-6.0055,-33.928,-27.393,-2.7965,-24.588,-3.0286,-33.792
827.0000000000,9053.8,982.57,1242.2,1507.0,1707.5,932.79,2702.9,326.22,1482.5,266.88,644.35,720.15,0.0000,-3728.8,-6748.2,-319.70,-2814.8,-2701.2,-13786.,-1697.6,-1354.9,-5245.0,-2893.1,-5711.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
828.0000000000,9060.7,969.44,1240.0,1502.5,1742.8,942.98,2692.1,326.05,1492.0,265.85,642.94,720.37,0.0000,-3765.6,-6765.1,-322.66,-2814.6,-2724.3,-13787.,-1697.6,-1373.4,-5254.2,-2894.3,-5717.4,2318.6,1036.4,793.89,745.09,1444.4,497.73,1784.1,515.56,788.16,235.26,338.11,407.27,0.0000,-2.4287,-2.5126,-0.37536,-2.2714,-1.6132,-9.1070,-7.3529,-0.75072,-6.6004,-0.81263,-9.0700
829.0000000000,9062.9,963.41,1240.6,1509.6,1746.8,937.37,2666.3,327.48,1498.6,267.12,640.49,723.48,0.0000,-3782.9,-6783.8,-325.55,-2814.6,-2732.2,-13787.,-1700.0,-1385.1,-5257.5,-2894.4,-5720.2,20435.,9134.1,6996.9,6566.9,12730.,4386.7,15724.,4543.9,6946.5,2073.4,2979.9,3589.5,0.0000,-21.444,-22.159,-3.3082,-20.038,-14.248,-80.260,-64.802,-6.6165,-58.172,-7.1606,-79.933
830.0000000000,9066.2,954.74,1234.5,1507.1,1693.8,918.10,2653.6,327.81,1487.7,264.73,648.75,729.82,0.0000,-3751.2,-6777.5,-323.79,-2814.5,-2710.2,-13785.,-1699.1,-1369.8,-5247.3,-2892.4,-5713.4,76.207,34.063,26.093,24.489,47.474,16.359,58.639,16.945,25.905,7.7324,11.113,13.386,0.0000,-0.79923E-01,-0.82643E-01,-0.12337E-01,-0.74667E-01,-0.53026E-01,-0.29929,-0.24165,-0.24674E-01,-0.21693,-0.26695E-01,-0.29806
831.0000000000,9071.9,946.37,1232.9,1496.9,1687.3,905.72,2654.5,330.21,1485.4,264.02,650.42,731.10,0.0000,-3740.0,-6767.7,-321.77,-2814.0,-2704.6,-13784.,-1698.2,-1362.8,-5244.1,-2891.7,-5710.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
832.0000000000,9066.8,946.79,1237.1,1496.6,1681.6,909.01,2656.7,331.37,1494.9,262.19,649.20,730.97,0.0000,-3777.3,-6781.8,-324.21,-2813.9,-2728.8,-13784.,-1699.5,-1381.7,-5254.7,-2893.8,-5718.4,14012.,6263.2,4797.8,4502.9,8729.0,3008.0,10782.,3115.7,4763.2,1421.7,2043.3,2461.3,0.0000,-14.705,-15.199,-2.2684,-13.735,-9.7588,-55.029,-44.426,-4.5369,-39.885,-4.9065,-54.795
833.0000000000,9069.4,943.93,1241.5,1501.2,1699.4,894.97,2664.2,333.75,1480.3,261.06,649.81,735.09,0.0000,-3793.8,-6798.4,-326.81,-2814.0,-2736.7,-13783.,-1708.9,-1392.9,-5259.7,-2894.5,-5723.4,76504.,34196.,26195.,24585.,47658.,16423.,58867.,17011.,26006.,7762.5,11156.,13438.,0.0000,-80.429,-83.036,-12.385,-75.061,-53.399,-300.46,-242.56,-24.770,-217.76,-26.786,-299.15
834.0000000000,9172.2,936.85,1242.0,1492.5,1692.3,875.98,2677.1,334.81,1480.0,259.64,647.58,732.17,0.0000,-3761.5,-6790.5,-324.87,-2813.9,-2714.6,-13782.,-1705.6,-1376.9,-5249.8,-2892.1,-5717.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
835.0000000000,9167.1,938.65,1231.4,1478.1,1682.2,868.86,2673.9,336.30,1474.2,258.48,641.64,732.55,0.0000,-3750.1,-6779.4,-322.71,-2813.6,-2708.8,-13781.,-1702.9,-1369.4,-5246.3,-2891.1,-5714.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
836.0000000000,9153.9,941.58,1252.6,1490.9,1687.6,883.44,2693.6,336.22,1476.9,260.20,641.44,736.65,0.0000,-3787.4,-6792.3,-325.06,-2813.4,-2733.0,-13781.,-1706.2,-1388.3,-5256.9,-2892.8,-5722.2,39737.,17762.,13606.,12770.,24754.,8530.2,30576.,8835.8,13508.,4031.9,5794.6,6979.9,0.0000,-41.779,-43.145,-6.4331,-38.972,-27.697,-156.09,-125.98,-12.866,-113.10,-13.904,-155.37
837.0000000000,9140.6,931.32,1245.3,1491.6,1708.0,902.12,2722.5,336.84,1464.9,263.88,642.33,736.07,0.0000,-3804.0,-6808.3,-327.58,-2813.9,-2741.3,-13781.,-1704.7,-1399.1,-5260.4,-2892.8,-5724.6,9608.8,4294.9,3290.0,3087.8,5985.9,2062.7,7393.6,2136.6,3266.3,974.96,1401.2,1687.8,0.0000,-10.121,-10.439,-1.5556,-9.4337,-6.7150,-37.750,-30.464,-3.1111,-27.348,-3.3615,-37.571
838.0000000000,9140.8,945.62,1245.1,1492.5,1722.9,920.12,2737.8,337.52,1468.4,264.25,642.27,726.81,0.0000,-3817.8,-6823.2,-329.68,-2814.6,-2747.7,-13782.,-1710.3,-1407.2,-5262.6,-2892.8,-5726.8,59357.,26531.,20324.,19075.,36977.,12742.,45673.,13198.,20177.,6022.7,8655.6,10426.,0.0000,-62.656,-64.534,-9.6094,-58.336,-41.588,-233.24,-188.21,-19.219,-168.95,-20.766,-232.11
839.0000000000,9144.1,957.42,1243.0,1484.8,1708.6,928.72,2746.3,333.01,1477.6,264.46,647.18,723.80,0.0000,-3830.7,-6836.8,-331.38,-2815.3,-2753.2,-13782.,-1706.7,-1413.9,-5263.0,-2892.7,-5727.2,1526.9,682.51,522.82,490.69,951.22,327.79,1174.9,339.53,519.05,154.93,222.66,268.21,0.0000,-1.6151,-1.6614,-0.24720,-1.5020,-1.0723,-6.0011,-4.8418,-0.49440,-4.3463,-0.53424,-5.9711
840.0000000000,9121.0,944.09,1236.8,1477.8,1655.3,905.90,2747.5,331.55,1464.9,265.30,647.69,720.64,0.0000,-3796.6,-6826.2,-328.68,-2815.3,-2729.9,-13782.,-1703.6,-1394.0,-5251.0,-2889.9,-5718.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
841.0000000000,9044.9,934.78,1248.2,1478.2,1653.0,909.91,2728.8,332.58,1462.4,268.80,646.45,726.12,0.0000,-3783.5,-6813.1,-325.98,-2815.3,-2724.3,-13781.,-1701.3,-1384.2,-5246.9,-2888.9,-5714.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
842.0000000000,9047.5,942.45,1241.9,1481.9,1644.7,911.86,2707.6,334.38,1467.7,266.19,647.75,728.89,0.0000,-3774.5,-6801.0,-323.86,-2814.9,-2720.0,-13782.,-1699.7,-1377.5,-5244.5,-2888.2,-5712.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
843.0000000000,9057.5,934.91,1242.1,1481.8,1643.9,902.35,2693.5,333.91,1460.0,264.39,643.92,728.06,0.0000,-3766.3,-6789.6,-322.23,-2814.6,-2716.4,-13782.,-1698.5,-1372.0,-5242.9,-2887.4,-5710.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
844.0000000000,8830.2,929.21,1240.5,1489.1,1652.8,913.15,2671.2,331.85,1471.1,267.05,643.14,733.69,0.0000,-3804.5,-6802.4,-325.05,-2814.9,-2741.0,-13783.,-1703.5,-1391.5,-5254.5,-2890.2,-5718.5,43332.,19369.,14837.,13925.,26994.,9302.0,33343.,9635.2,14730.,4396.7,6318.8,7611.4,0.0000,-45.739,-47.119,-7.0151,-42.564,-30.340,-170.40,-137.43,-14.030,-123.36,-15.147,-169.50
845.0000000000,8680.6,917.55,1225.6,1489.8,1679.3,907.68,2658.8,328.98,1464.0,264.85,642.57,737.58,0.0000,-3775.6,-6793.9,-323.82,-2815.1,-2720.7,-13783.,-1701.4,-1377.7,-5246.2,-2888.7,-5713.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
846.0000000000,8695.4,909.05,1224.2,1487.0,1669.8,896.43,2657.4,331.07,1464.8,265.24,639.91,734.61,0.0000,-3764.7,-6782.8,-322.26,-2814.7,-2715.1,-13783.,-1699.8,-1370.8,-5243.2,-2887.9,-5710.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
847.0000000000,8681.4,901.35,1227.2,1498.8,1668.8,899.39,2655.6,333.14,1479.5,265.95,638.39,734.96,0.0000,-3801.9,-6795.5,-325.02,-2814.1,-2738.9,-13783.,-1708.3,-1390.0,-5255.0,-2889.8,-5720.1,72767.,32525.,24915.,23384.,45331.,15621.,55992.,16180.,24736.,7383.3,10611.,12782.,0.0000,-76.756,-79.094,-11.780,-71.463,-50.872,-286.10,-230.79,-23.561,-207.15,-25.417,-284.59
848.0000000000,8681.7,898.22,1213.5,1495.4,1680.2,871.83,2674.7,330.86,1459.0,262.96,637.86,732.93,0.0000,-3772.6,-6787.4,-323.75,-2813.3,-2718.1,-13782.,-1705.0,-1376.4,-5246.8,-2887.8,-5715.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
849.0000000000,8675.1,915.39,1205.0,1493.6,1686.4,864.86,2697.8,328.24,1439.9,262.86,635.85,730.78,0.0000,-3761.7,-6777.5,-322.17,-2812.4,-2712.4,-13782.,-1702.3,-1369.8,-5243.6,-2886.8,-5712.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
850.0000000000,8733.2,917.27,1188.6,1493.2,1687.3,876.94,2734.2,328.97,1441.5,266.21,639.02,735.41,0.0000,-3753.7,-6767.6,-320.86,-2811.8,-2708.9,-13782.,-1700.3,-1365.2,-5241.6,-2886.1,-5711.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
851.0000000000,8799.5,932.10,1180.9,1490.1,1666.1,882.80,2732.0,332.28,1449.5,266.54,646.59,734.42,0.0000,-3747.6,-6758.8,-319.82,-2811.3,-2706.1,-13782.,-1698.8,-1361.5,-5240.3,-2885.8,-5709.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
852.0000000000,8831.3,905.64,1213.0,1492.3,1649.4,864.68,2708.8,333.81,1444.7,269.39,645.32,733.73,0.0000,-3741.3,-6751.3,-318.98,-2810.6,-2702.9,-13782.,-1697.8,-1358.1,-5239.5,-2885.5,-5708.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
853.0000000000,8842.6,909.64,1213.8,1501.7,1646.9,865.55,2706.0,334.28,1437.0,267.93,645.67,734.05,0.0000,-3735.3,-6744.2,-318.27,-2810.0,-2699.9,-13782.,-1697.0,-1355.1,-5238.6,-2885.2,-5707.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
854.0000000000,8853.1,913.56,1219.5,1517.5,1652.6,874.38,2717.0,337.99,1443.2,266.66,646.98,735.98,0.0000,-3729.9,-6737.7,-317.66,-2809.5,-2696.9,-13781.,-1696.4,-1352.6,-5238.0,-2885.2,-5706.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
855.0000000000,8839.3,903.38,1224.4,1518.0,1656.2,881.55,2729.5,337.30,1447.8,264.67,648.33,737.77,0.0000,-3724.4,-6732.6,-317.10,-2808.9,-2693.7,-13780.,-1696.1,-1350.2,-5237.3,-2884.7,-5706.0,613.94,274.42,210.21,197.29,382.46,131.79,472.40,136.51,208.70,62.293,89.526,107.84,0.0000,-0.64282,-0.66524,-0.99391E-01,-0.60090,-0.42470,-2.4145,-1.9471,-0.19878,-1.7477,-0.21410,-2.4009
856.0000000000,8843.3,903.57,1200.0,1508.6,1652.3,877.40,2729.8,336.74,1443.2,262.98,645.03,735.90,0.0000,-3719.1,-6727.6,-316.59,-2808.2,-2690.8,-13779.,-1695.8,-1348.0,-5236.6,-2884.1,-5705.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
857.0000000000,8839.9,902.88,1177.4,1513.0,1655.5,894.55,2696.1,337.77,1441.6,260.15,640.08,736.38,0.0000,-3759.4,-6745.3,-320.18,-2808.0,-2716.0,-13779.,-1695.8,-1368.7,-5247.3,-2886.3,-5713.0,1705.3,762.23,583.89,548.00,1062.3,366.07,1312.2,379.18,579.68,173.03,248.67,299.53,0.0000,-1.7863,-1.8472,-0.27607,-1.6706,-1.1811,-6.7059,-5.4078,-0.55214,-4.8543,-0.59438,-6.6676
858.0000000000,8852.2,894.41,1177.4,1509.9,1649.6,892.79,2682.2,338.51,1434.9,259.94,638.57,733.20,0.0000,-3732.9,-6742.3,-319.54,-2807.6,-2696.3,-13778.,-1695.6,-1358.1,-5239.0,-2884.5,-5707.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
859.0000000000,8847.7,894.02,1179.1,1511.9,1642.9,887.86,2678.0,337.34,1439.9,260.80,638.53,736.52,0.0000,-3724.3,-6735.6,-318.41,-2807.0,-2691.4,-13777.,-1695.4,-1353.3,-5236.4,-2883.6,-5706.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
860.0000000000,8824.9,891.02,1176.8,1505.1,1638.4,869.54,2683.3,338.67,1450.4,259.85,640.56,735.23,0.0000,-3717.9,-6729.0,-317.41,-2806.3,-2688.1,-13776.,-1695.2,-1350.1,-5235.2,-2883.0,-5705.2,1.6564,0.74040,0.56717,0.53231,1.0319,0.35559,1.2746,0.36832,0.56308,0.16807,0.24155,0.29096,0.0000,-0.17311E-02,-0.17928E-02,-0.26816E-03,-0.16205E-02,-0.11418E-02,-0.65133E-02,-0.52521E-02,-0.53633E-03,-0.47149E-02,-0.57692E-03,-0.64751E-02
861.0000000000,8811.5,899.64,1185.8,1506.3,1651.8,882.58,2690.8,337.92,1437.6,259.82,639.47,734.50,0.0000,-3757.4,-6746.7,-320.67,-2806.0,-2713.2,-13776.,-1725.3,-1370.2,-5252.3,-2885.5,-5720.7,0.22588E+06,0.10096E+06,77340.,72586.,0.14071E+06,48489.,0.17381E+06,50225.,76783.,22919.,32938.,39676.,0.0000,-236.42,-244.52,-36.567,-221.25,-156.13,-888.15,-716.34,-73.135,-642.94,-78.659,-882.94
862.0000000000,8804.0,914.93,1188.1,1482.7,1648.5,888.79,2697.1,340.48,1434.8,261.90,634.68,740.70,0.0000,-3776.3,-6766.7,-323.87,-2805.8,-2721.6,-13777.,-1740.1,-1382.8,-5263.0,-2886.2,-5733.1,0.16639E+06,74372.,56971.,53469.,0.10365E+06,35718.,0.12803E+06,36997.,56560.,16882.,24263.,29226.,0.0000,-174.50,-180.23,-26.937,-163.16,-115.27,-654.32,-527.82,-53.873,-473.62,-57.933,-650.48
863.0000000000,8810.2,1018.5,1242.7,1490.0,1650.2,995.97,2818.4,354.35,1431.5,279.40,664.77,783.19,0.0000,-3796.1,-6787.5,-326.52,-2807.6,-2733.4,-13781.,-1744.8,-1392.3,-5270.5,-2888.8,-5741.7,0.12221E+06,54626.,41845.,39273.,76131.,26234.,94037.,27174.,41543.,12400.,17821.,21466.,0.0000,-128.79,-132.59,-19.785,-120.19,-85.438,-481.45,-388.02,-39.569,-348.05,-42.641,-478.30
864.0000000000,8818.6,1063.6,1286.5,1506.4,1632.7,991.14,2817.6,350.31,1429.0,297.22,682.38,793.63,0.0000,-3815.7,-6808.8,-328.67,-2809.8,-2741.9,-13787.,-1737.6,-1400.4,-5277.3,-2892.5,-5744.9,46515.,20791.,15927.,14948.,28977.,9985.3,35792.,10343.,15812.,4719.7,6783.0,8170.5,0.0000,-49.206,-50.523,-7.5304,-45.835,-32.722,-183.45,-147.79,-15.061,-132.53,-16.257,-182.20
865.0000000000,8817.6,1110.9,1291.9,1512.9,1621.5,961.64,2775.8,356.24,1424.4,294.96,701.74,823.98,0.0000,-3833.2,-6824.8,-330.45,-2812.6,-2747.9,-13791.,-1729.1,-1407.5,-5279.4,-2897.0,-5745.2,24814.,11091.,8496.3,7974.0,15458.,5326.7,19093.,5517.5,8435.0,2517.7,3618.4,4358.6,0.0000,-26.316,-26.973,-4.0171,-24.480,-17.514,-97.899,-78.873,-8.0343,-70.715,-8.6789,-97.239
866.0000000000,8836.9,1110.7,1308.0,1515.2,1575.2,931.52,2748.8,367.41,1428.7,285.51,726.53,807.57,0.0000,-3846.9,-6840.5,-332.07,-2813.7,-2752.4,-13793.,-1732.2,-1414.5,-5280.8,-2902.3,-5746.5,93821.,41936.,32124.,30150.,58446.,20140.,72192.,20862.,31893.,9519.6,13681.,16480.,0.0000,-99.653,-102.05,-15.189,-92.613,-66.293,-370.09,-298.31,-30.378,-267.40,-32.812,-367.75
867.0000000000,8855.7,1127.6,1302.4,1511.4,1604.9,925.49,2770.6,376.36,1437.7,285.44,754.88,806.55,0.0000,-3859.3,-6855.2,-333.52,-2813.8,-2757.3,-13796.,-1744.7,-1421.1,-5284.2,-2908.2,-5751.6,0.16733E+06,74795.,57295.,53774.,0.10424E+06,35921.,0.12876E+06,37208.,56882.,16979.,24401.,29393.,0.0000,-178.03,-182.16,-27.090,-165.28,-118.37,-660.05,-532.26,-54.180,-476.98,-58.520,-656.10
868.0000000000,8867.3,1191.2,1423.5,1508.4,1604.1,1012.4,2934.0,396.76,1422.1,306.57,762.94,840.70,0.0000,-3830.7,-6846.1,-330.76,-2814.8,-2737.9,-13802.,-1731.5,-1401.2,-5274.0,-2910.2,-5744.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
869.0000000000,8892.4,1240.3,1458.2,1514.4,1622.1,978.07,2946.5,396.18,1432.2,317.92,770.02,861.62,0.0000,-3823.7,-6832.6,-328.14,-2816.5,-2731.9,-13807.,-1721.6,-1391.6,-5272.1,-2913.7,-5739.5,865.10,386.68,296.21,278.00,538.92,185.71,665.67,192.36,294.07,87.777,126.15,151.96,0.0000,-0.92180,-0.94260,-0.14005,-0.85465,-0.61330,-3.4183,-2.7546,-0.28010,-2.4676,-0.30332,-3.3973
870.0000000000,8906.5,1269.5,1529.9,1515.6,1652.5,937.12,2911.1,403.64,1458.7,313.72,809.33,851.04,0.0000,-3817.1,-6824.1,-326.23,-2816.3,-2726.6,-13811.,-1714.3,-1385.5,-5269.0,-2919.0,-5736.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
871.0000000000,8902.5,1259.1,1526.1,1514.7,1719.3,977.95,2940.3,417.81,1472.7,312.78,793.23,833.70,0.0000,-3858.7,-6836.2,-328.93,-2815.8,-2749.9,-13816.,-1719.0,-1405.2,-5278.7,-2923.1,-5744.6,73321.,32773.,25105.,23562.,45676.,15740.,56418.,16303.,24924.,7439.5,10692.,12879.,0.0000,-78.087,-79.877,-11.870,-72.431,-51.905,-289.50,-233.51,-23.740,-209.16,-25.686,-288.00
872.0000000000,8920.6,1246.5,1561.3,1525.9,1722.4,982.31,2987.9,402.04,1473.7,323.38,765.41,836.46,0.0000,-3877.2,-6850.6,-331.74,-2815.6,-2756.4,-13819.,-1715.0,-1416.1,-5281.9,-2923.9,-5747.9,15168.,6780.0,5193.6,4874.4,9449.2,3256.2,11672.,3372.8,5156.2,1539.1,2211.9,2664.4,0.0000,-16.173,-16.534,-2.4556,-14.993,-10.749,-59.866,-48.309,-4.9112,-43.271,-5.3095,-59.575
873.0000000000,8949.7,1194.5,1594.0,1534.9,1773.7,997.71,2942.0,398.79,1484.3,326.90,753.01,848.79,0.0000,-3891.6,-6864.9,-334.02,-2816.3,-2761.1,-13820.,-1710.6,-1424.4,-5282.3,-2923.9,-5749.6,3983.8,1780.7,1364.1,1280.2,2481.8,855.20,3065.4,885.83,1354.2,404.22,580.94,699.77,0.0000,-4.2543,-4.3466,-0.64495,-3.9405,-2.8276,-15.720,-12.688,-1.2899,-11.365,-1.3939,-15.645
874.0000000000,8972.0,1187.7,1655.7,1541.2,1830.8,992.23,2973.4,395.96,1516.1,332.81,738.91,864.90,0.0000,-3905.4,-6879.7,-335.85,-2817.3,-2766.1,-13823.,-1712.6,-1432.8,-5283.9,-2922.9,-5751.6,43409.,19403.,14863.,13950.,27042.,9318.5,33402.,9652.3,14756.,4404.5,6330.0,7624.8,0.0000,-46.443,-47.411,-7.0275,-42.972,-30.871,-171.28,-138.25,-14.055,-123.84,-15.184,-170.46
875.0000000000,8977.7,1179.9,1659.7,1564.1,1934.5,1056.4,2949.4,385.64,1543.4,344.18,748.10,836.43,0.0000,-3918.5,-6892.8,-337.33,-2821.1,-2771.7,-13826.,-1709.0,-1439.1,-5286.5,-2922.6,-5751.7,4004.2,1789.8,1371.0,1286.7,2494.4,859.56,3081.1,890.35,1361.1,406.28,583.90,703.34,0.0000,-4.2937,-4.3779,-0.64824,-3.9675,-2.8551,-15.801,-12.753,-1.2965,-11.424,-1.4005,-15.724
876.0000000000,9004.8,1184.5,1639.5,1567.2,1861.1,1056.0,2905.2,381.24,1553.9,336.93,733.90,829.10,0.0000,-3931.0,-6907.4,-338.55,-2824.4,-2776.6,-13828.,-1708.2,-1444.5,-5286.4,-2921.8,-5751.2,18248.,8156.5,6248.1,5864.1,11368.,3917.3,14041.,4057.6,6203.1,1851.5,2661.0,3205.3,0.0000,-19.610,-19.971,-2.9542,-18.094,-13.039,-72.014,-58.120,-5.9084,-52.061,-6.3813,-71.660
877.0000000000,9004.2,1147.3,1607.1,1571.5,1876.7,1088.3,2905.3,380.01,1555.7,339.70,714.92,820.41,0.0000,-3896.3,-6895.2,-335.46,-2829.0,-2754.7,-13829.,-1705.2,-1423.0,-5274.0,-2917.4,-5742.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
878.0000000000,9029.5,1139.2,1611.7,1580.3,1901.3,1116.6,2872.9,373.40,1570.6,339.86,723.39,805.58,0.0000,-3883.3,-6877.8,-332.50,-2833.2,-2749.3,-13831.,-1703.0,-1411.5,-5269.1,-2914.9,-5737.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
879.0000000000,9046.1,1153.9,1600.7,1576.0,1870.4,1096.8,2872.8,370.40,1549.9,334.29,721.50,799.89,0.0000,-3919.0,-6885.5,-334.31,-2836.2,-2773.2,-13834.,-1726.8,-1428.9,-5282.2,-2915.9,-5750.4,0.18923E+06,84582.,64792.,60810.,0.11788E+06,40621.,0.14561E+06,42077.,64325.,19200.,27594.,33238.,0.0000,-203.34,-207.24,-30.635,-187.60,-135.24,-746.88,-602.80,-61.269,-539.87,-66.118,-743.13
880.0000000000,9033.1,1149.4,1576.2,1578.3,1901.8,1107.0,2901.4,370.50,1544.7,336.17,723.86,809.49,0.0000,-3933.3,-6895.2,-336.46,-2838.8,-2781.3,-13837.,-1719.9,-1438.1,-5286.2,-2916.3,-5755.4,3298.7,1474.5,1129.5,1060.1,2055.0,708.13,2538.3,733.50,1121.3,334.71,481.03,579.43,0.0000,-3.5516,-3.6156,-0.53404,-3.2746,-2.3656,-13.025,-10.510,-1.0681,-9.4120,-1.1525,-12.959
881.0000000000,8903.1,1206.7,1602.9,1577.2,1878.0,1136.2,2949.2,382.64,1540.7,340.77,760.25,826.93,0.0000,-3948.4,-6907.8,-338.36,-2841.5,-2788.7,-13843.,-1733.7,-1444.8,-5291.8,-2918.2,-5761.4,0.14716E+06,65778.,50388.,47291.,91675.,31591.,0.11324E+06,32722.,50025.,14932.,21460.,25849.,0.0000,-159.08,-161.55,-23.824,-146.37,-106.14,-581.56,-469.09,-47.648,-419.98,-51.511,-578.33
882.0000000000,8904.3,1129.0,1608.6,1577.4,1846.5,1122.1,2895.3,395.66,1559.5,340.89,753.90,833.70,0.0000,-3913.5,-6896.3,-335.80,-2844.1,-2765.6,-13846.,-1724.1,-1424.0,-5282.4,-2917.0,-5754.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
883.0000000000,8972.6,1130.7,1642.4,1581.6,1915.7,1130.7,2932.9,406.74,1563.2,350.72,809.74,848.65,0.0000,-3902.3,-6887.1,-333.29,-2846.7,-2760.8,-13850.,-1716.7,-1413.9,-5279.6,-2919.6,-5750.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
884.0000000000,8959.0,1168.7,1630.6,1593.3,1908.2,1061.0,2881.4,402.73,1559.0,354.00,820.20,864.25,0.0000,-3893.0,-6875.3,-331.39,-2848.9,-2756.0,-13852.,-1711.2,-1406.9,-5278.4,-2923.4,-5747.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
885.0000000000,8954.3,1156.5,1628.7,1600.9,1912.1,1051.2,2884.7,425.64,1566.9,357.20,819.13,858.32,0.0000,-3885.0,-6864.5,-330.01,-2850.0,-2751.8,-13854.,-1707.3,-1401.3,-5275.9,-2926.6,-5745.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
886.0000000000,8950.2,1132.5,1641.0,1601.1,1895.5,1061.4,2945.6,428.76,1577.7,350.35,796.80,822.10,0.0000,-3878.0,-6852.5,-328.98,-2850.2,-2747.2,-13856.,-1704.7,-1396.5,-5273.1,-2926.9,-5742.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
887.0000000000,8903.0,1163.3,1588.4,1607.8,1901.1,1085.5,2979.8,413.91,1598.4,353.13,765.66,829.21,0.0000,-3871.3,-6839.1,-328.16,-2850.5,-2742.9,-13857.,-1702.8,-1391.7,-5271.4,-2925.2,-5741.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
888.0000000000,8918.0,1153.3,1628.6,1614.3,1908.7,1078.5,2968.3,402.43,1600.0,356.52,742.57,828.14,0.0000,-3865.0,-6828.7,-327.48,-2850.9,-2738.8,-13858.,-1701.5,-1387.4,-5269.4,-2922.4,-5740.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
889.0000000000,8903.5,1149.9,1627.5,1626.9,1960.5,1073.1,2959.0,405.66,1609.8,354.00,745.36,828.17,0.0000,-3857.8,-6819.8,-326.91,-2850.7,-2735.1,-13862.,-1700.6,-1383.8,-5267.4,-2920.4,-5740.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
890.0000000000,8905.0,1101.8,1632.3,1627.9,1941.9,1077.2,2952.6,404.65,1603.4,355.04,751.31,834.13,0.0000,-3850.1,-6812.9,-326.40,-2850.7,-2731.7,-13864.,-1699.9,-1380.6,-5266.1,-2920.9,-5740.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
891.0000000000,8922.9,1085.1,1626.2,1634.3,1894.3,1085.2,2986.8,409.17,1627.1,356.00,744.19,845.44,0.0000,-3842.8,-6805.6,-325.90,-2851.1,-2728.6,-13866.,-1699.5,-1379.0,-5265.5,-2921.0,-5740.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
892.0000000000,8945.8,1079.3,1648.7,1644.3,1911.0,1089.2,3018.3,405.58,1615.8,356.48,733.65,837.72,0.0000,-3837.3,-6798.9,-325.41,-2851.2,-2725.1,-13868.,-1699.2,-1377.7,-5265.7,-2919.1,-5740.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
893.0000000000,8942.0,1114.0,1622.6,1663.8,1929.1,1134.0,3035.7,400.84,1626.2,358.59,731.55,819.69,0.0000,-3831.6,-6791.7,-324.93,-2852.6,-2721.8,-13870.,-1698.9,-1375.4,-5266.2,-2916.6,-5740.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
894.0000000000,8953.5,1132.3,1624.6,1668.5,1855.9,1153.0,3018.9,395.18,1674.1,358.27,715.38,825.34,0.0000,-3872.0,-6811.3,-328.55,-2853.5,-2746.7,-13871.,-1700.9,-1396.8,-5277.0,-2917.0,-5748.4,15416.,6890.6,5278.4,4954.0,9603.4,3309.3,11862.,3427.8,5240.3,1564.2,2248.0,2707.8,0.0000,-16.463,-16.864,-2.4957,-15.289,-11.009,-60.901,-49.130,-4.9914,-43.999,-5.4034,-60.572
895.0000000000,9011.2,1084.6,1622.3,1685.4,1854.6,1184.0,2994.7,396.91,1676.4,358.78,709.10,827.73,0.0000,-3889.9,-6832.6,-331.97,-2855.8,-2755.8,-13872.,-1717.1,-1409.7,-5283.4,-2916.9,-5755.8,0.12475E+06,55759.,42713.,40088.,77712.,26779.,95988.,27738.,42405.,12657.,18191.,21912.,0.0000,-133.43,-136.53,-20.195,-123.85,-89.313,-492.76,-397.58,-40.391,-356.03,-43.724,-490.10
896.0000000000,9044.5,1063.8,1632.1,1715.2,1860.8,1194.0,3001.0,396.93,1690.9,358.47,718.48,823.57,0.0000,-3904.2,-6850.6,-334.68,-2857.1,-2762.0,-13872.,-1714.3,-1419.4,-5286.4,-2917.2,-5759.6,13799.,6167.9,4724.8,4434.4,8596.2,2962.2,10618.,3068.3,4690.7,1400.1,2012.2,2423.8,0.0000,-14.787,-15.113,-2.2339,-13.712,-9.9022,-54.503,-43.978,-4.4679,-39.382,-4.8368,-54.208
897.0000000000,9043.4,1079.1,1614.2,1745.8,1869.2,1191.8,3005.9,389.79,1666.1,356.58,715.03,816.33,0.0000,-3916.8,-6866.7,-336.80,-2858.6,-2767.3,-13872.,-1718.1,-1427.8,-5288.1,-2917.2,-5762.9,59396.,26549.,20337.,19087.,37001.,12750.,45703.,13207.,20190.,6026.6,8661.3,10433.,0.0000,-63.772,-65.104,-9.6156,-59.072,-42.711,-234.60,-189.30,-19.231,-169.51,-20.820,-233.32
898.0000000000,9050.0,1112.0,1595.5,1772.1,1903.1,1187.5,3006.8,388.11,1655.1,356.46,717.75,820.87,0.0000,-3928.2,-6880.5,-338.48,-2860.6,-2772.8,-13872.,-1716.3,-1435.4,-5288.9,-2917.1,-5764.4,25004.,11176.,8561.3,8035.1,15576.,5367.5,19240.,5559.8,8499.6,2537.0,3646.2,4392.0,0.0000,-26.899,-27.431,-4.0479,-24.891,-18.027,-98.773,-79.692,-8.0958,-71.359,-8.7657,-98.229
899.0000000000,9046.8,1143.2,1575.6,1792.3,1863.2,1207.6,3023.9,393.06,1639.9,354.61,722.21,817.20,0.0000,-3939.7,-6890.7,-339.88,-2862.8,-2778.5,-13873.,-1711.9,-1442.2,-5288.2,-2917.4,-5764.1,3470.4,1551.2,1188.3,1115.2,2161.9,744.98,2670.3,771.66,1179.7,352.12,506.06,609.58,0.0000,-3.7425,-3.8108,-0.56182,-3.4581,-2.5097,-13.713,-11.061,-1.1236,-9.9046,-1.2172,-13.635
900.0000000000,9123.0,1135.1,1590.6,1796.0,1850.8,1237.2,3062.8,401.80,1642.1,357.33,726.40,812.90,0.0000,-3951.4,-6902.5,-341.08,-2864.8,-2784.0,-13875.,-1708.4,-1448.4,-5287.0,-2917.8,-5762.8,1359.6,607.71,465.52,436.91,846.97,291.86,1046.2,302.32,462.17,137.95,198.26,238.82,0.0000,-1.4700,-1.4951,-0.22011,-1.3561,-0.98626,-5.3744,-4.3338,-0.44021,-3.8806,-0.47722,-5.3424
901.0000000000,9163.2,1118.8,1584.1,1795.1,1853.6,1237.4,3078.3,402.37,1661.3,356.68,724.24,798.69,0.0000,-3961.5,-6914.1,-342.13,-2866.3,-2788.4,-13876.,-1713.5,-1454.1,-5287.9,-2917.4,-5763.2,57840.,25853.,19804.,18587.,36032.,12416.,44506.,12861.,19662.,5868.8,8434.4,10160.,0.0000,-62.648,-63.675,-9.3638,-57.730,-42.041,-228.66,-184.38,-18.728,-165.09,-20.305,-227.28
902.0000000000,9176.6,1132.4,1571.2,1798.2,1862.4,1258.6,3086.1,394.56,1649.7,348.53,722.25,788.20,0.0000,-3970.8,-6923.0,-343.05,-2867.6,-2792.5,-13876.,-1710.5,-1459.2,-5287.4,-2916.5,-5762.7,6129.2,2739.6,2098.6,1969.6,3818.2,1315.7,4716.2,1362.9,2083.5,621.90,893.78,1076.6,0.0000,-6.6493,-6.7547,-0.99226,-6.1212,-4.4630,-24.232,-19.539,-1.9845,-17.495,-2.1517,-24.085
903.0000000000,9184.7,1132.0,1529.1,1787.7,1870.6,1268.2,3095.9,390.29,1634.2,348.95,728.26,784.55,0.0000,-3932.7,-6907.4,-339.76,-2868.8,-2768.2,-13876.,-1707.2,-1436.6,-5275.3,-2913.8,-5753.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
904.0000000000,9219.2,1141.4,1517.2,1794.4,1856.9,1279.8,3072.1,395.66,1637.0,349.64,733.94,788.55,0.0000,-3962.7,-6914.4,-340.74,-2870.0,-2788.9,-13876.,-1706.9,-1451.7,-5282.6,-2915.0,-5758.1,14563.,6509.3,4986.3,4679.8,9072.0,3126.2,11206.,3238.1,4950.3,1477.6,2123.6,2558.0,0.0000,-15.796,-16.056,-2.3576,-14.539,-10.599,-57.576,-46.423,-4.7152,-41.566,-5.1120,-57.224
905.0000000000,9276.6,1141.1,1515.3,1777.4,1838.6,1258.9,3087.9,403.07,1612.7,345.32,731.09,786.88,0.0000,-3928.1,-6900.9,-338.07,-2870.2,-2766.9,-13875.,-1704.8,-1432.5,-5271.4,-2912.7,-5750.6,745.61,333.27,255.29,239.60,464.48,160.06,573.72,165.79,253.45,75.653,108.73,130.97,0.0000,-0.80784,-0.82189,-0.12071,-0.74375,-0.54174,-2.9482,-2.3768,-0.24141,-2.1282,-0.26179,-2.9298
906.0000000000,9177.4,1132.1,1511.1,1779.4,1823.5,1243.9,3094.2,413.75,1596.0,342.72,732.03,791.22,0.0000,-3912.9,-6885.8,-335.49,-2870.1,-2760.2,-13875.,-1703.1,-1422.6,-5267.6,-2911.8,-5747.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
907.0000000000,8998.0,1109.5,1511.6,1764.4,1805.1,1248.3,3050.2,412.01,1607.3,339.67,727.73,792.17,0.0000,-3900.6,-6870.7,-333.45,-2869.8,-2755.3,-13872.,-1701.9,-1415.4,-5265.6,-2911.4,-5744.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
908.0000000000,8930.5,1129.7,1527.2,1779.4,1799.1,1254.7,3071.6,422.40,1634.5,337.98,731.25,795.60,0.0000,-3936.2,-6880.1,-335.96,-2869.6,-2779.1,-13871.,-1711.1,-1435.1,-5277.6,-2913.8,-5754.0,74292.,33207.,25437.,23874.,46281.,15948.,57165.,16519.,25254.,7538.0,10833.,13049.,0.0000,-80.325,-81.805,-12.027,-74.069,-53.912,-293.73,-236.81,-24.054,-212.04,-26.089,-291.85
909.0000000000,8909.3,1153.6,1534.0,1781.1,1797.5,1227.0,3085.9,430.77,1614.7,333.84,734.01,791.63,0.0000,-3951.0,-6893.5,-338.58,-2869.5,-2785.8,-13870.,-1717.2,-1444.9,-5282.7,-2914.7,-5759.4,67430.,30140.,23088.,21669.,42006.,14475.,51885.,14993.,22921.,6841.7,9832.8,11844.,0.0000,-73.012,-74.301,-10.916,-67.281,-49.018,-266.59,-214.94,-21.832,-192.45,-23.683,-264.87
910.0000000000,8886.8,1144.9,1528.3,1768.8,1784.1,1217.6,3056.5,432.06,1616.7,337.13,725.99,783.74,0.0000,-3962.1,-6906.4,-340.69,-2869.4,-2790.5,-13871.,-1713.0,-1451.9,-5283.9,-2914.6,-5761.2,3611.0,1614.0,1236.4,1160.4,2249.5,775.16,2778.5,802.93,1227.5,366.39,526.57,634.28,0.0000,-3.9155,-3.9824,-0.58459,-3.6053,-2.6288,-14.276,-11.510,-1.1692,-10.306,-1.2683,-14.184
911.0000000000,8899.0,1131.7,1523.2,1765.9,1792.9,1225.6,3071.3,433.45,1597.1,341.77,724.02,782.12,0.0000,-3925.7,-6894.1,-338.24,-2869.4,-2767.7,-13870.,-1709.2,-1431.5,-5271.9,-2912.1,-5752.8,313.95,140.33,107.50,100.89,195.58,67.396,241.58,69.810,106.72,31.855,45.782,55.147,0.0000,-0.34009,-0.34627,-0.50826E-01,-0.31326,-0.22830,-1.2416,-1.0008,-0.10165,-0.89607,-0.11029,-1.2334
912.0000000000,8898.9,1147.8,1536.7,1776.7,1770.7,1263.5,3071.2,433.79,1608.5,344.76,736.58,789.16,0.0000,-3958.8,-6904.3,-339.81,-2869.6,-2789.5,-13871.,-1708.7,-1447.7,-5279.5,-2914.2,-5757.3,17525.,7833.3,6000.5,5631.7,10917.,3762.0,13485.,3896.8,5957.2,1778.2,2555.5,3078.3,0.0000,-19.026,-19.344,-2.8371,-17.506,-12.783,-69.327,-55.870,-5.6742,-50.022,-6.1623,-68.854
913.0000000000,8863.4,1150.5,1534.5,1766.7,1773.4,1251.3,3065.1,432.39,1608.1,345.47,731.10,786.36,0.0000,-3925.2,-6892.3,-337.53,-2869.4,-2767.2,-13871.,-1706.0,-1429.4,-5269.9,-2912.0,-5749.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
914.0000000000,8686.4,1136.7,1556.3,1729.4,1798.4,1266.6,3076.4,432.67,1616.9,347.85,727.62,791.53,0.0000,-3911.0,-6877.6,-335.18,-2868.9,-2760.1,-13870.,-1704.0,-1419.9,-5266.3,-2911.3,-5746.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
915.0000000000,8682.9,1114.8,1568.6,1713.1,1834.5,1256.2,3088.6,430.34,1649.1,347.21,723.76,790.79,0.0000,-3899.9,-6864.0,-333.27,-2867.7,-2754.7,-13869.,-1702.6,-1412.9,-5264.0,-2910.3,-5744.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
916.0000000000,8669.5,1103.4,1596.0,1717.4,1822.8,1251.5,3062.5,424.15,1651.9,351.64,713.91,789.53,0.0000,-3889.5,-6851.6,-331.77,-2866.3,-2750.0,-13869.,-1701.6,-1407.1,-5262.5,-2909.7,-5743.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
917.0000000000,8686.8,1121.0,1615.0,1749.8,1804.3,1260.4,3043.4,419.59,1670.0,350.39,720.63,788.34,0.0000,-3880.0,-6840.7,-330.57,-2865.4,-2745.9,-13871.,-1700.8,-1402.4,-5261.1,-2909.6,-5742.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
918.0000000000,8723.4,1130.0,1600.4,1760.0,1798.3,1252.6,3020.6,424.29,1695.2,348.52,725.17,787.49,0.0000,-3871.2,-6831.3,-329.55,-2864.6,-2742.2,-13872.,-1700.4,-1398.5,-5259.6,-2909.9,-5741.5,507.09,226.66,173.63,162.95,315.89,108.86,390.19,112.75,172.37,51.452,73.945,89.071,0.0000,-0.54529,-0.55751,-0.82093E-01,-0.50415,-0.36582,-2.0037,-1.6161,-0.16419,-1.4472,-0.17820,-1.9913
919.0000000000,8741.5,1130.4,1605.6,1755.5,1788.2,1266.4,3015.9,426.63,1732.4,344.29,720.03,783.90,0.0000,-3909.6,-6846.4,-332.76,-2864.1,-2766.6,-13874.,-1710.3,-1419.8,-5271.6,-2912.3,-5751.7,75945.,33946.,26003.,24405.,47310.,16303.,58437.,16887.,25816.,7705.8,11075.,13340.,0.0000,-81.784,-83.498,-12.295,-75.581,-54.914,-300.01,-242.04,-24.590,-216.73,-26.688,-298.20
920.0000000000,8728.2,1115.7,1565.8,1753.2,1745.2,1267.0,3048.7,419.03,1729.7,337.94,710.98,781.55,0.0000,-3879.8,-6838.7,-331.79,-2863.4,-2745.9,-13875.,-1707.5,-1406.6,-5263.2,-2910.0,-5747.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
921.0000000000,8766.5,1102.5,1557.6,1767.0,1736.2,1280.6,3067.2,416.31,1727.7,336.03,708.57,777.66,0.0000,-3868.0,-6828.3,-330.41,-2862.7,-2740.2,-13877.,-1705.1,-1400.5,-5259.8,-2908.9,-5745.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
922.0000000000,8781.6,1088.4,1544.0,1757.0,1745.6,1276.5,3056.0,417.48,1718.7,338.14,712.64,773.59,0.0000,-3858.9,-6818.1,-329.18,-2862.1,-2735.9,-13878.,-1703.4,-1396.3,-5258.1,-2907.9,-5744.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
923.0000000000,8818.9,1094.9,1537.2,1758.8,1733.8,1269.4,3035.1,415.16,1688.5,337.34,714.74,774.45,0.0000,-3851.0,-6810.8,-328.14,-2861.6,-2732.1,-13879.,-1702.0,-1392.8,-5256.6,-2906.9,-5743.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
924.0000000000,8827.7,1093.8,1511.4,1777.1,1755.6,1298.2,3003.7,411.35,1681.7,338.78,701.28,773.74,0.0000,-3843.7,-6804.1,-327.26,-2861.4,-2728.9,-13878.,-1701.1,-1389.6,-5255.4,-2905.8,-5742.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
925.0000000000,8823.5,1105.0,1514.8,1786.9,1729.2,1317.7,2988.8,413.70,1695.0,334.96,696.44,776.25,0.0000,-3837.2,-6797.7,-326.50,-2861.2,-2726.1,-13877.,-1700.4,-1386.7,-5254.4,-2904.8,-5741.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
926.0000000000,8822.5,1111.3,1529.5,1793.2,1713.0,1323.7,2999.6,411.54,1699.4,329.14,693.39,776.36,0.0000,-3830.7,-6792.2,-325.82,-2860.8,-2723.2,-13876.,-1699.9,-1384.0,-5253.6,-2904.2,-5740.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
927.0000000000,8811.0,1102.2,1533.3,1784.0,1705.4,1289.4,3029.5,417.49,1688.7,334.14,686.33,776.75,0.0000,-3824.0,-6787.4,-325.19,-2860.4,-2720.3,-13874.,-1699.6,-1381.0,-5253.2,-2903.3,-5740.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
928.0000000000,8805.1,1093.0,1534.6,1772.5,1736.0,1266.6,3017.3,413.89,1674.6,338.04,680.40,787.50,0.0000,-3817.6,-6781.9,-324.60,-2860.4,-2717.7,-13873.,-1699.3,-1378.7,-5252.7,-2902.8,-5739.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
929.0000000000,8787.8,1098.9,1534.3,1779.6,1744.5,1248.3,2979.7,412.78,1650.4,336.43,686.22,796.87,0.0000,-3811.8,-6776.7,-324.04,-2860.3,-2715.1,-13871.,-1699.1,-1376.4,-5251.9,-2902.5,-5739.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
930.0000000000,8652.1,1096.6,1527.6,1781.5,1733.8,1252.7,2941.4,415.33,1641.2,336.58,684.48,791.89,0.0000,-3806.0,-6771.3,-323.52,-2860.2,-2712.5,-13868.,-1699.0,-1374.3,-5251.2,-2902.2,-5738.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
931.0000000000,8602.2,1096.8,1499.2,1778.4,1737.8,1228.0,2929.1,420.10,1671.0,335.41,686.42,791.89,0.0000,-3800.1,-6765.6,-323.01,-2859.8,-2710.0,-13865.,-1698.8,-1372.3,-5250.5,-2901.6,-5738.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
932.0000000000,8601.3,1086.0,1506.9,1762.5,1725.0,1218.7,2915.6,418.17,1675.3,333.14,688.30,780.42,0.0000,-3794.5,-6760.2,-322.54,-2859.3,-2707.6,-13863.,-1698.7,-1370.4,-5250.0,-2901.3,-5737.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
933.0000000000,8598.9,1097.5,1509.2,1742.5,1662.9,1227.8,2957.2,416.97,1670.3,331.90,693.37,784.46,0.0000,-3789.1,-6756.0,-322.08,-2858.2,-2705.1,-13862.,-1698.6,-1368.5,-5249.5,-2901.1,-5737.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
934.0000000000,8557.0,1076.9,1534.0,1750.2,1582.7,1246.3,2939.7,415.17,1668.1,333.01,688.57,784.09,0.0000,-3784.0,-6752.8,-321.58,-2857.1,-2702.7,-13859.,-1698.5,-1366.6,-5249.1,-2900.6,-5737.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
935.0000000000,8533.9,1079.2,1519.3,1745.7,1525.3,1245.5,2955.6,406.05,1697.7,336.47,681.44,782.56,0.0000,-3779.0,-6749.2,-321.07,-2856.1,-2700.4,-13857.,-1698.5,-1364.9,-5248.7,-2899.9,-5737.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
936.0000000000,8506.5,1090.8,1530.7,1749.2,1540.6,1263.3,2987.9,412.11,1706.0,339.33,679.26,782.95,0.0000,-3774.2,-6746.0,-320.55,-2855.1,-2698.1,-13855.,-1698.4,-1363.5,-5248.0,-2899.2,-5736.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
937.0000000000,8507.1,1074.2,1544.0,1727.2,1545.2,1243.0,2989.4,409.44,1736.6,335.67,680.03,785.82,0.0000,-3769.7,-6743.3,-320.05,-2854.1,-2695.8,-13853.,-1698.3,-1362.2,-5247.6,-2898.3,-5736.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
938.0000000000,8459.8,1072.4,1561.4,1735.7,1572.4,1236.9,2986.9,414.29,1750.5,335.92,675.66,785.67,0.0000,-3765.1,-6740.2,-319.60,-2853.1,-2693.6,-13852.,-1698.2,-1360.6,-5247.2,-2897.2,-5736.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
939.0000000000,8465.0,1057.5,1575.6,1753.6,1600.4,1286.6,2968.1,412.50,1801.2,336.65,683.31,782.32,0.0000,-3760.3,-6735.9,-319.18,-2852.1,-2691.4,-13850.,-1698.1,-1359.2,-5246.7,-2896.2,-5735.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
940.0000000000,8495.5,1108.5,1570.6,1752.3,1558.9,1283.7,2930.0,408.84,1848.8,334.70,688.96,783.35,0.0000,-3755.6,-6732.0,-318.76,-2851.0,-2689.1,-13848.,-1698.0,-1357.9,-5246.2,-2895.4,-5735.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
941.0000000000,8690.1,1133.2,1550.1,1758.9,1535.2,1250.3,2913.1,410.71,1842.5,342.74,687.62,791.61,0.0000,-3750.8,-6728.6,-318.35,-2849.7,-2686.8,-13847.,-1698.0,-1356.6,-5245.7,-2894.6,-5735.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
942.0000000000,8846.5,1175.7,1556.0,1775.2,1539.1,1251.2,2908.3,413.73,1827.9,344.25,677.17,795.28,0.0000,-3745.9,-6725.3,-317.96,-2848.4,-2684.4,-13844.,-1697.9,-1355.4,-5245.2,-2893.9,-5734.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
943.0000000000,8860.6,1207.8,1586.5,1794.9,1542.2,1275.3,2916.5,408.19,1822.7,348.69,664.29,798.68,0.0000,-3786.3,-6745.1,-321.64,-2847.5,-2710.1,-13843.,-1700.7,-1376.4,-5257.1,-2895.9,-5743.4,21042.,9405.2,7204.6,6761.8,13108.,4516.9,16191.,4678.7,7152.7,2135.0,3068.3,3696.0,0.0000,-22.156,-22.862,-3.4064,-20.758,-14.803,-82.918,-66.937,-6.8129,-59.979,-7.3705,-82.387
944.0000000000,8856.0,1184.7,1592.1,1795.5,1539.6,1293.6,2931.4,407.29,1844.4,350.79,656.29,801.63,0.0000,-3805.2,-6766.8,-325.13,-2846.9,-2719.1,-13841.,-1702.8,-1390.0,-5261.2,-2896.4,-5747.0,21371.,9552.3,7317.3,6867.6,13313.,4587.6,16444.,4751.9,7264.6,2168.4,3116.3,3753.8,0.0000,-22.544,-23.231,-3.4597,-21.104,-15.068,-84.201,-67.980,-6.9195,-60.915,-7.4863,-83.666
945.0000000000,8881.3,1166.6,1592.3,1775.7,1550.5,1283.5,2934.8,406.03,1866.2,345.55,653.76,800.18,0.0000,-3774.6,-6763.5,-323.82,-2845.9,-2697.6,-13839.,-1701.5,-1376.5,-5251.3,-2894.0,-5740.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
946.0000000000,8895.4,1160.7,1615.1,1766.0,1562.1,1247.7,2919.1,406.31,1886.4,339.99,654.55,795.15,0.0000,-3763.9,-6755.8,-322.11,-2844.8,-2692.4,-13836.,-1700.3,-1370.6,-5248.3,-2893.0,-5737.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
947.0000000000,8715.3,1145.6,1599.9,1755.6,1503.3,1232.2,2939.7,403.75,1882.2,335.41,648.37,788.24,0.0000,-3756.1,-6748.3,-320.69,-2843.7,-2689.1,-13834.,-1699.5,-1366.7,-5246.8,-2892.2,-5736.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
948.0000000000,8702.4,1129.4,1587.5,1747.0,1474.1,1223.4,2949.4,401.16,1850.3,327.41,648.12,792.43,0.0000,-3749.3,-6741.7,-319.56,-2842.6,-2686.4,-13833.,-1698.8,-1363.6,-5245.7,-2891.6,-5735.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
949.0000000000,8637.9,1097.7,1578.2,1748.3,1476.3,1213.4,2969.6,408.59,1792.0,321.95,639.84,791.33,0.0000,-3743.1,-6735.8,-318.65,-2841.6,-2684.0,-13832.,-1698.3,-1361.2,-5244.8,-2891.0,-5734.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
950.0000000000,8477.5,1050.6,1583.7,1755.6,1468.6,1253.7,3006.7,419.48,1780.2,321.38,635.39,773.49,0.0000,-3737.5,-6729.9,-317.91,-2840.6,-2681.7,-13831.,-1697.9,-1359.1,-5243.9,-2890.0,-5733.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
951.0000000000,8333.6,1054.4,1551.0,1759.2,1472.8,1250.7,3042.6,422.57,1761.9,319.69,632.43,773.57,0.0000,-3732.1,-6724.0,-317.27,-2839.6,-2679.5,-13830.,-1697.6,-1357.3,-5243.4,-2889.1,-5733.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
952.0000000000,8326.7,1076.5,1546.4,1770.6,1504.0,1243.3,3054.1,416.87,1791.8,321.68,629.00,767.84,0.0000,-3726.9,-6718.5,-316.71,-2838.8,-2677.4,-13828.,-1697.4,-1355.5,-5243.0,-2888.3,-5732.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
953.0000000000,8349.2,1079.9,1566.7,1791.7,1511.9,1255.4,3047.3,416.49,1789.3,327.31,631.56,767.55,0.0000,-3722.0,-6713.4,-316.22,-2837.9,-2675.5,-13825.,-1697.2,-1353.6,-5242.6,-2887.5,-5731.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
954.0000000000,8392.4,1112.0,1557.7,1789.6,1564.3,1273.4,3063.5,412.44,1792.7,332.10,637.95,771.27,0.0000,-3717.5,-6708.9,-315.73,-2837.0,-2673.5,-13823.,-1697.1,-1351.7,-5242.3,-2886.8,-5731.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
955.0000000000,8310.1,1164.3,1551.4,1791.2,1582.2,1323.3,3025.6,409.32,1804.3,342.29,637.78,777.99,0.0000,-3758.0,-6727.9,-319.31,-2836.4,-2699.6,-13821.,-1699.9,-1372.1,-5254.0,-2888.8,-5739.3,21211.,9480.8,7262.6,6816.2,13213.,4553.3,16321.,4716.4,7210.2,2152.2,3093.0,3725.7,0.0000,-22.226,-22.979,-3.4338,-20.869,-14.774,-83.458,-67.409,-6.8677,-60.428,-7.4201,-82.932
956.0000000000,8171.2,1179.4,1670.6,1814.4,1543.9,1328.3,3022.9,405.17,1827.5,345.44,632.23,777.73,0.0000,-3777.3,-6748.7,-322.71,-2836.0,-2708.7,-13819.,-1701.3,-1385.1,-5257.8,-2889.3,-5742.4,15953.,7130.9,5462.5,5126.7,9938.3,3424.7,12276.,3547.4,5423.1,1618.7,2326.4,2802.3,0.0000,-16.749,-17.291,-2.5827,-15.713,-11.138,-62.768,-50.698,-5.1654,-45.449,-5.5808,-62.371
957.0000000000,8073.5,1178.4,1687.0,1817.7,1527.2,1317.4,3024.4,397.20,1859.8,344.02,625.92,788.46,0.0000,-3793.0,-6767.9,-325.41,-2835.6,-2715.8,-13817.,-1704.4,-1395.3,-5259.8,-2889.6,-5744.4,32168.,14379.,11014.,10337.,20039.,6905.5,24752.,7152.8,10935.,3263.9,4690.9,5650.4,0.0000,-33.840,-34.886,-5.2077,-31.711,-22.502,-126.56,-102.22,-10.415,-91.639,-11.252,-125.75
958.0000000000,7855.5,1138.9,1668.3,1805.3,1534.1,1338.3,3038.4,396.99,1895.4,342.07,623.20,785.53,0.0000,-3807.1,-6785.0,-327.52,-2835.4,-2721.9,-13814.,-1708.7,-1404.0,-5262.0,-2889.7,-5746.5,46352.,20718.,15871.,14895.,28875.,9950.3,35666.,10307.,15756.,4703.1,6759.2,8141.8,0.0000,-48.857,-50.302,-7.5040,-45.728,-32.481,-182.36,-147.30,-15.008,-132.04,-16.212,-181.19
959.0000000000,7844.3,1121.5,1677.2,1800.3,1526.8,1327.7,2997.1,392.36,1877.7,339.16,623.45,782.12,0.0000,-3773.9,-6776.6,-325.11,-2834.8,-2699.5,-13812.,-1705.5,-1386.9,-5251.1,-2887.1,-5738.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
960.0000000000,7712.8,1106.1,1699.8,1799.9,1589.0,1344.5,3002.3,391.75,1872.2,333.69,628.72,770.00,0.0000,-3761.5,-6764.5,-322.61,-2834.0,-2693.8,-13810.,-1702.9,-1378.8,-5247.1,-2885.8,-5735.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
961.0000000000,7665.0,1097.8,1710.1,1790.4,1595.6,1326.5,3001.2,392.20,1870.9,332.33,632.31,767.09,0.0000,-3752.3,-6752.8,-320.61,-2833.1,-2690.1,-13808.,-1701.0,-1373.4,-5244.9,-2884.8,-5733.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
962.0000000000,7648.1,1107.6,1712.2,1788.9,1599.1,1341.4,3004.1,401.79,1870.4,332.42,631.84,764.34,0.0000,-3790.1,-6765.8,-323.15,-2832.4,-2715.5,-13808.,-1708.2,-1392.8,-5256.8,-2886.6,-5741.6,64148.,28673.,21964.,20614.,39961.,13770.,49359.,14264.,21806.,6508.7,9354.2,11268.,0.0000,-67.557,-69.608,-10.385,-63.213,-44.820,-252.43,-203.83,-20.770,-182.72,-22.419,-250.73
963.0000000000,7656.6,1122.2,1746.8,1788.1,1617.9,1369.3,3011.2,406.34,1836.3,331.72,642.06,759.65,0.0000,-3807.6,-6781.8,-325.83,-2831.7,-2724.1,-13808.,-1709.0,-1404.0,-5260.8,-2887.3,-5744.9,28142.,12579.,9635.7,9043.4,17531.,6041.1,21654.,6257.5,9566.2,2855.4,4103.7,4943.1,0.0000,-29.699,-30.554,-4.5559,-27.761,-19.717,-110.77,-89.428,-9.1118,-80.164,-9.8376,-110.00
964.0000000000,7426.0,1107.6,1756.9,1788.0,1616.5,1319.4,3072.1,404.72,1817.8,333.57,647.44,750.59,0.0000,-3775.5,-6774.6,-323.93,-2830.7,-2702.2,-13807.,-1705.5,-1387.4,-5250.5,-2884.6,-5737.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
965.0000000000,7307.5,1115.1,1730.5,1772.2,1575.3,1274.2,3100.9,404.30,1809.1,336.92,642.66,751.18,0.0000,-3763.6,-6763.5,-321.78,-2829.6,-2696.5,-13806.,-1702.9,-1379.5,-5247.1,-2883.2,-5734.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
966.0000000000,7223.3,1118.3,1729.2,1751.5,1535.3,1292.9,3108.8,405.08,1789.1,333.72,640.43,755.72,0.0000,-3754.9,-6753.0,-320.02,-2828.6,-2693.3,-13804.,-1700.9,-1374.0,-5245.3,-2882.2,-5731.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
967.0000000000,7193.4,1156.2,1746.2,1739.3,1500.4,1310.4,3107.7,411.76,1762.0,333.53,651.88,757.88,0.0000,-3748.0,-6744.6,-318.65,-2827.7,-2690.7,-13803.,-1699.5,-1369.6,-5244.0,-2881.6,-5729.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
968.0000000000,7192.5,1155.9,1725.0,1752.1,1475.0,1302.6,3063.4,408.39,1790.9,333.45,648.68,759.16,0.0000,-3786.9,-6760.4,-321.62,-2827.0,-2716.2,-13803.,-1700.2,-1389.5,-5255.2,-2883.7,-5735.5,12242.,5472.1,4191.8,3934.1,7626.4,2628.0,9420.1,2722.2,4161.5,1242.2,1785.2,2150.4,0.0000,-12.897,-13.284,-1.9819,-12.059,-8.5490,-48.213,-38.905,-3.9638,-34.876,-4.2775,-47.857
969.0000000000,7164.6,1143.0,1710.7,1788.2,1499.9,1321.1,3031.2,417.51,1781.6,331.64,639.63,760.96,0.0000,-3804.6,-6778.3,-324.59,-2826.7,-2724.7,-13801.,-1701.2,-1400.9,-5258.5,-2884.5,-5737.3,15420.,6892.2,5279.6,4955.1,9605.7,3310.1,11865.,3428.6,5241.6,1564.5,2248.5,2708.5,0.0000,-16.270,-16.740,-2.4963,-15.202,-10.789,-60.724,-49.002,-4.9926,-43.927,-5.3869,-60.277
970.0000000000,7127.6,1134.1,1688.9,1784.6,1486.9,1288.9,3050.1,418.47,1763.5,328.61,634.85,768.94,0.0000,-3772.8,-6770.7,-322.89,-2826.3,-2702.9,-13799.,-1699.8,-1384.5,-5248.0,-2882.4,-5729.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
971.0000000000,7107.6,1080.6,1703.2,1784.9,1529.3,1288.1,3053.7,425.71,1723.4,329.08,631.95,769.92,0.0000,-3761.2,-6759.7,-320.88,-2825.4,-2697.1,-13797.,-1698.7,-1376.7,-5244.6,-2881.2,-5726.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
972.0000000000,7097.8,1018.8,1717.3,1762.2,1527.6,1302.0,3064.5,425.67,1705.0,330.20,625.36,769.04,0.0000,-3752.2,-6749.2,-319.22,-2824.3,-2693.3,-13796.,-1697.8,-1371.3,-5243.0,-2880.1,-5724.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
973.0000000000,7097.5,994.36,1740.8,1767.1,1583.0,1297.4,3077.2,427.15,1658.1,325.45,620.22,760.64,0.0000,-3790.0,-6763.1,-321.99,-2823.4,-2717.9,-13795.,-1698.4,-1390.6,-5253.7,-2882.1,-5731.3,8317.2,3717.6,2847.8,2672.8,5181.2,1785.4,6399.8,1849.4,2827.3,843.90,1212.8,1460.9,0.0000,-8.7620,-9.0250,-1.3465,-8.1894,-5.7945,-32.751,-26.426,-2.6929,-23.692,-2.9026,-32.505
974.0000000000,7111.8,1018.6,1722.6,1756.6,1598.4,1260.8,3085.3,421.37,1661.2,322.93,619.36,749.05,0.0000,-3761.1,-6756.4,-320.76,-2822.5,-2697.8,-13793.,-1697.6,-1377.4,-5245.0,-2880.2,-5725.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
975.0000000000,7118.0,1027.0,1712.3,1756.1,1572.4,1227.9,3079.6,422.02,1657.2,325.87,620.34,743.56,0.0000,-3750.4,-6746.5,-319.20,-2821.4,-2692.6,-13792.,-1697.0,-1370.8,-5242.3,-2879.5,-5722.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
976.0000000000,7106.6,1013.8,1700.3,1752.1,1550.5,1244.0,3092.3,417.30,1638.1,327.68,622.59,744.48,0.0000,-3742.2,-6736.9,-317.89,-2820.2,-2688.9,-13790.,-1696.6,-1366.1,-5240.8,-2878.8,-5721.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
977.0000000000,7137.5,1037.7,1684.7,1739.7,1540.3,1244.7,3086.4,415.46,1643.3,324.46,623.62,743.27,0.0000,-3735.0,-6728.1,-316.83,-2818.8,-2685.7,-13789.,-1696.2,-1362.3,-5239.7,-2878.3,-5720.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
978.0000000000,7168.5,1041.0,1696.9,1728.1,1517.1,1220.1,3066.8,415.43,1667.5,322.29,621.96,741.13,0.0000,-3728.3,-6720.2,-315.96,-2817.3,-2682.7,-13789.,-1695.9,-1359.0,-5238.8,-2878.0,-5719.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
979.0000000000,7190.5,1085.9,1679.5,1722.8,1523.1,1222.7,3078.0,410.21,1711.5,323.87,618.32,741.51,0.0000,-3721.9,-6713.4,-315.21,-2815.8,-2680.0,-13788.,-1695.7,-1356.1,-5238.0,-2877.7,-5718.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
980.0000000000,7200.8,1123.7,1665.5,1716.5,1524.2,1220.9,3071.7,404.96,1687.7,322.51,613.76,758.57,0.0000,-3716.3,-6707.5,-314.55,-2814.4,-2677.3,-13787.,-1695.5,-1353.5,-5237.4,-2877.4,-5718.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
981.0000000000,7125.8,1101.5,1665.6,1719.1,1518.8,1222.3,3055.1,404.17,1688.2,321.88,617.50,753.18,0.0000,-3711.1,-6702.1,-313.97,-2813.0,-2674.8,-13786.,-1695.3,-1351.2,-5236.9,-2877.1,-5717.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
982.0000000000,7133.0,1109.7,1681.2,1708.7,1517.9,1225.5,3047.2,410.84,1657.1,322.32,612.97,752.72,0.0000,-3706.1,-6697.2,-313.43,-2811.7,-2672.2,-13784.,-1695.2,-1349.2,-5236.4,-2876.7,-5717.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
983.0000000000,7147.6,1130.5,1710.7,1720.6,1510.5,1242.4,3008.6,416.94,1663.5,318.79,613.50,745.63,0.0000,-3746.3,-6715.8,-316.98,-2810.7,-2697.6,-13784.,-1700.1,-1369.8,-5248.4,-2878.6,-5726.5,37197.,16626.,12736.,11953.,23172.,7985.0,28622.,8271.1,12644.,3774.2,5424.2,6533.7,0.0000,-38.895,-40.211,-6.0219,-36.491,-25.581,-146.50,-118.11,-12.044,-105.92,-12.945,-145.24
984.0000000000,7156.5,1121.8,1697.7,1701.1,1509.0,1208.8,3023.7,420.98,1651.3,315.88,609.20,740.45,0.0000,-3719.8,-6712.8,-316.31,-2809.6,-2678.2,-13783.,-1698.8,-1359.5,-5240.3,-2876.5,-5721.5,145.21,64.904,49.718,46.662,90.457,31.171,111.73,32.288,49.360,14.733,21.174,25.506,0.0000,-0.15174,-0.15694,-0.23508E-01,-0.14236,-0.99661E-01,-0.57188,-0.46105,-0.47015E-01,-0.41347,-0.50516E-01,-0.56694
985.0000000000,7166.4,1139.9,1710.7,1672.1,1507.1,1225.1,2996.4,423.40,1654.5,315.24,607.72,740.42,0.0000,-3756.3,-6729.7,-319.22,-2808.8,-2701.5,-13782.,-1700.6,-1377.8,-5249.8,-2878.1,-5728.5,21783.,9736.6,7458.5,7000.0,13570.,4676.1,16761.,4843.6,7404.7,2210.2,3176.5,3826.2,0.0000,-22.800,-23.549,-3.5265,-21.378,-14.985,-85.787,-69.162,-7.0529,-62.025,-7.5767,-85.042
986.0000000000,7179.4,1148.8,1732.4,1659.9,1499.2,1219.1,2995.1,419.98,1613.0,315.67,602.90,735.84,0.0000,-3728.1,-6724.8,-317.99,-2807.7,-2681.3,-13781.,-1699.0,-1365.7,-5240.9,-2875.8,-5722.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
987.0000000000,7215.0,1154.1,1727.9,1658.2,1488.2,1223.0,2982.1,418.54,1619.4,313.72,600.78,730.60,0.0000,-3718.5,-6716.7,-316.41,-2806.5,-2676.2,-13780.,-1697.7,-1360.0,-5237.8,-2874.6,-5720.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
988.0000000000,7152.2,1161.9,1704.0,1646.0,1474.1,1202.8,2986.8,417.32,1617.7,316.11,600.14,737.02,0.0000,-3711.5,-6708.6,-315.08,-2805.3,-2672.7,-13779.,-1696.7,-1356.2,-5236.3,-2873.8,-5719.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
989.0000000000,7033.8,1168.9,1693.9,1656.5,1422.1,1192.9,2976.0,414.91,1612.0,318.85,592.70,734.37,0.0000,-3705.3,-6701.2,-314.01,-2804.0,-2669.5,-13777.,-1696.0,-1353.2,-5235.2,-2873.1,-5718.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
990.0000000000,7001.2,1175.8,1693.8,1647.1,1420.3,1182.9,2968.4,414.56,1616.6,315.15,593.53,734.72,0.0000,-3699.6,-6694.5,-313.13,-2802.9,-2666.6,-13775.,-1695.5,-1350.6,-5234.5,-2872.5,-5717.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
991.0000000000,6975.0,1189.4,1697.0,1626.7,1405.9,1184.8,2976.8,412.18,1616.1,312.84,586.68,734.78,0.0000,-3694.2,-6688.5,-312.43,-2801.9,-2663.8,-13773.,-1695.1,-1348.2,-5233.9,-2871.9,-5716.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
992.0000000000,6960.5,1188.7,1689.7,1626.7,1410.3,1199.0,2987.9,413.17,1624.5,312.85,588.16,735.32,0.0000,-3689.0,-6683.1,-311.82,-2800.9,-2661.3,-13772.,-1694.8,-1346.0,-5233.4,-2871.3,-5715.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
993.0000000000,6997.1,1167.2,1697.6,1625.2,1425.6,1203.3,3030.7,415.00,1609.4,318.59,593.88,735.63,0.0000,-3684.0,-6678.1,-311.30,-2800.1,-2658.9,-13770.,-1694.5,-1343.9,-5233.1,-2870.7,-5715.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
994.0000000000,7004.2,1160.4,1708.2,1627.0,1435.8,1199.1,3069.4,416.48,1597.5,320.68,595.46,741.80,0.0000,-3679.3,-6673.4,-310.82,-2799.1,-2656.7,-13769.,-1694.3,-1342.1,-5232.7,-2870.1,-5715.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
995.0000000000,7017.1,1142.9,1710.4,1621.5,1433.0,1205.4,3059.0,420.20,1588.3,318.27,594.85,748.83,0.0000,-3674.9,-6668.8,-310.38,-2798.2,-2654.4,-13767.,-1694.2,-1340.4,-5232.3,-2869.5,-5714.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
996.0000000000,7046.5,1144.9,1709.7,1600.5,1424.9,1222.6,3053.5,417.79,1590.2,316.60,594.97,745.32,0.0000,-3670.4,-6665.0,-309.95,-2797.3,-2652.1,-13766.,-1694.0,-1338.8,-5231.9,-2868.8,-5714.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
997.0000000000,7029.9,1122.7,1717.3,1593.9,1416.4,1222.3,3037.2,415.42,1584.0,315.96,596.69,736.50,0.0000,-3666.2,-6661.3,-309.55,-2796.4,-2649.9,-13764.,-1693.9,-1337.3,-5231.5,-2868.2,-5714.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
998.0000000000,6797.4,1130.9,1694.4,1571.5,1439.1,1206.6,3016.1,412.94,1585.8,318.37,607.08,739.30,0.0000,-3662.1,-6658.1,-309.16,-2795.5,-2647.6,-13763.,-1693.7,-1335.8,-5231.3,-2867.6,-5713.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
999.0000000000,6805.7,1144.4,1681.1,1563.4,1473.9,1197.3,2996.6,415.36,1566.1,321.71,610.54,731.92,0.0000,-3658.0,-6655.4,-308.78,-2794.6,-2645.5,-13761.,-1693.6,-1334.4,-5231.0,-2866.9,-5713.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1000.000000000,6796.0,1133.3,1672.1,1567.3,1467.6,1217.6,2978.3,419.37,1556.0,326.07,616.33,735.90,0.0000,-3698.7,-6675.7,-312.45,-2793.9,-2671.3,-13760.,-1695.6,-1354.6,-5242.6,-2868.8,-5721.7,15269.,6824.8,5228.0,4906.6,9511.7,3277.7,11749.,3395.1,5190.3,1549.2,2226.5,2682.0,0.0000,-15.818,-16.411,-2.4719,-14.902,-10.318,-60.081,-48.436,-4.9437,-43.455,-5.3025,-59.533
1001.000000000,6662.7,1114.6,1683.0,1569.7,1475.3,1224.5,2977.0,422.93,1533.1,326.17,614.28,733.43,0.0000,-3673.1,-6674.2,-311.90,-2793.0,-2652.3,-13758.,-1695.0,-1345.4,-5234.6,-2866.7,-5716.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1002.000000000,6562.4,1133.4,1738.8,1566.2,1467.6,1202.2,2990.1,424.34,1533.6,323.35,613.37,728.77,0.0000,-3665.3,-6669.2,-310.82,-2791.8,-2647.9,-13757.,-1694.5,-1341.2,-5232.3,-2865.7,-5714.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1003.000000000,6523.6,1110.3,1727.7,1548.3,1467.1,1187.3,3003.1,427.78,1532.6,323.49,616.02,725.07,0.0000,-3659.7,-6663.9,-309.87,-2790.6,-2645.1,-13755.,-1694.1,-1338.4,-5231.4,-2864.9,-5713.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1004.000000000,6430.3,1109.3,1705.9,1539.2,1481.6,1191.3,2996.9,432.26,1529.0,322.67,621.58,729.83,0.0000,-3654.5,-6659.0,-309.08,-2789.5,-2642.6,-13753.,-1693.7,-1336.2,-5230.8,-2864.2,-5713.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1005.000000000,6384.2,1109.4,1703.7,1536.5,1500.6,1193.9,2985.6,439.26,1524.9,322.96,629.77,730.29,0.0000,-3649.8,-6654.5,-308.42,-2788.3,-2640.4,-13751.,-1693.4,-1334.2,-5230.4,-2863.5,-5712.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1006.000000000,6362.1,1080.8,1700.0,1526.5,1512.5,1187.5,2988.5,441.33,1521.2,324.59,635.40,728.48,0.0000,-3645.2,-6650.4,-307.86,-2787.2,-2638.3,-13749.,-1693.2,-1332.4,-5229.9,-2862.9,-5711.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1007.000000000,6377.0,1075.9,1690.9,1501.2,1503.2,1179.1,2966.7,449.60,1499.0,324.92,636.75,730.78,0.0000,-3640.8,-6646.8,-307.35,-2786.1,-2636.2,-13747.,-1693.1,-1330.7,-5229.4,-2862.0,-5711.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1008.000000000,6376.9,1073.4,1690.1,1497.8,1608.5,1162.6,2983.4,452.14,1496.9,325.84,636.16,723.46,0.0000,-3636.4,-6643.5,-306.87,-2785.0,-2634.2,-13745.,-1692.9,-1329.1,-5228.8,-2861.3,-5711.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1009.000000000,6371.9,1072.6,1730.9,1500.0,1848.6,1142.7,2972.3,456.21,1483.2,324.85,633.45,726.56,0.0000,-3632.1,-6640.3,-306.41,-2784.0,-2632.2,-13743.,-1692.8,-1327.7,-5228.4,-2860.8,-5710.7,444.97,198.89,152.36,142.99,277.20,95.521,342.39,98.943,151.26,45.149,64.887,78.160,0.0000,-0.45786,-0.47668,-0.72037E-01,-0.43277,-0.29682,-1.7507,-1.4107,-0.14407,-1.2660,-0.15443,-1.7333
1010.000000000,6381.0,1070.9,1742.0,1512.0,1841.4,1140.4,2929.9,457.74,1491.9,321.85,628.75,724.33,0.0000,-3628.0,-6637.4,-305.98,-2782.9,-2630.2,-13741.,-1692.7,-1326.5,-5227.8,-2860.2,-5710.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1011.000000000,6390.3,1056.6,1743.1,1524.4,1853.4,1126.8,2897.3,460.14,1516.7,322.38,625.98,727.79,0.0000,-3624.3,-6634.4,-305.56,-2781.9,-2628.3,-13740.,-1692.6,-1325.7,-5227.3,-2859.7,-5709.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1012.000000000,6438.1,1070.8,1758.1,1541.7,1858.2,1142.6,2863.4,456.94,1537.1,323.64,617.10,727.43,0.0000,-3665.1,-6654.3,-309.17,-2781.0,-2654.4,-13739.,-1715.9,-1345.7,-5243.1,-2861.7,-5723.5,0.17473E+06,78100.,59826.,56149.,0.10885E+06,37508.,0.13445E+06,38852.,59395.,17729.,25479.,30691.,0.0000,-179.84,-187.06,-28.287,-169.92,-116.62,-687.40,-553.93,-56.573,-497.08,-60.633,-680.44
1013.000000000,6444.6,1079.6,1776.0,1507.6,1858.5,1134.1,2855.8,451.00,1556.9,327.32,614.93,731.27,0.0000,-3684.6,-6676.5,-312.63,-2780.3,-2663.6,-13739.,-1713.6,-1359.2,-5249.2,-2862.2,-5729.9,27265.,12187.,9335.5,8761.7,16985.,5852.9,20980.,6062.6,9268.2,2766.5,3975.9,4789.2,0.0000,-28.123,-29.206,-4.4140,-26.546,-18.242,-107.26,-86.441,-8.8279,-77.566,-9.4615,-106.17
1014.000000000,6449.9,1097.7,1783.6,1500.7,1856.3,1109.6,2854.6,448.98,1538.2,325.72,615.84,735.93,0.0000,-3655.7,-6673.8,-311.32,-2779.5,-2642.8,-13737.,-1707.8,-1347.1,-5239.0,-2859.7,-5723.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1015.000000000,6406.9,1120.3,1819.0,1500.1,1869.7,1137.1,2864.0,455.21,1556.2,329.16,620.43,733.83,0.0000,-3647.6,-6667.4,-309.64,-2779.1,-2639.2,-13737.,-1703.3,-1341.6,-5235.0,-2859.2,-5720.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1016.000000000,6367.1,1120.6,1833.0,1498.7,1861.9,1143.6,2838.2,458.98,1560.7,330.86,624.76,738.88,0.0000,-3642.2,-6662.1,-308.25,-2778.4,-2636.5,-13738.,-1700.0,-1338.1,-5232.4,-2858.6,-5717.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1017.000000000,6211.0,1133.3,1821.6,1472.1,1821.4,1146.1,2838.7,456.87,1574.8,333.30,620.09,736.39,0.0000,-3637.3,-6656.8,-307.17,-2777.5,-2634.0,-13738.,-1697.6,-1335.4,-5230.9,-2858.2,-5715.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1018.000000000,6217.1,1117.7,1822.2,1466.9,1818.2,1143.2,2855.7,454.23,1593.3,334.09,621.93,729.23,0.0000,-3632.6,-6651.8,-306.30,-2776.5,-2631.6,-13737.,-1696.0,-1333.1,-5229.6,-2857.7,-5713.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1019.000000000,6236.8,1156.8,1788.6,1448.1,1826.8,1121.7,2846.9,448.58,1604.7,332.32,620.95,736.21,0.0000,-3628.2,-6647.2,-305.58,-2775.7,-2629.0,-13736.,-1694.8,-1331.1,-5228.5,-2857.4,-5712.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1020.000000000,6226.3,1145.3,1765.4,1442.2,1835.3,1131.2,2829.2,444.83,1609.0,330.63,623.43,738.18,0.0000,-3624.0,-6642.7,-304.99,-2774.8,-2626.7,-13736.,-1694.0,-1329.3,-5227.5,-2857.0,-5710.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1021.000000000,6146.8,1131.4,1763.6,1440.0,1840.1,1147.1,2828.2,443.06,1609.6,328.22,620.79,741.71,0.0000,-3619.8,-6638.8,-304.48,-2773.7,-2624.4,-13735.,-1693.3,-1327.7,-5226.4,-2856.4,-5709.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1022.000000000,6077.0,1126.9,1780.6,1443.8,1841.6,1158.6,2841.5,442.28,1587.0,328.27,617.43,737.01,0.0000,-3615.7,-6635.3,-304.03,-2772.4,-2622.2,-13735.,-1692.9,-1326.2,-5225.3,-2855.7,-5709.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1023.000000000,6116.4,1138.2,1788.8,1450.8,1831.0,1157.9,2839.4,442.91,1601.2,326.84,624.45,726.37,0.0000,-3611.9,-6631.9,-303.62,-2771.2,-2620.1,-13734.,-1692.5,-1324.8,-5224.6,-2855.4,-5708.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1024.000000000,6334.2,1158.8,1804.5,1449.0,1820.1,1136.3,2847.5,436.52,1598.9,321.88,626.26,728.69,0.0000,-3608.1,-6629.7,-303.27,-2770.0,-2618.1,-13734.,-1692.3,-1323.6,-5223.9,-2855.1,-5708.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1025.000000000,6475.6,1170.5,1779.2,1443.7,1604.0,1145.5,2839.0,443.92,1631.9,320.42,628.87,728.57,0.0000,-3648.8,-6650.4,-306.95,-2768.9,-2644.1,-13735.,-1693.5,-1343.1,-5235.0,-2857.3,-5716.0,10812.,4832.9,3702.1,3474.6,6735.6,2321.0,8319.7,2404.2,3675.4,1097.1,1576.7,1899.2,0.0000,-11.094,-11.548,-1.7504,-10.496,-7.1558,-42.545,-34.280,-3.5008,-30.763,-3.7505,-42.106
1026.000000000,6470.8,1189.3,1769.0,1448.7,1509.3,1172.5,2838.8,445.08,1611.9,320.51,631.18,726.20,0.0000,-3668.4,-6673.0,-310.48,-2768.1,-2653.4,-13735.,-1695.6,-1356.2,-5238.6,-2858.1,-5719.3,19138.,8554.2,6552.8,6150.0,11922.,4108.3,14726.,4255.4,6505.5,1941.8,2790.7,3361.6,0.0000,-19.678,-20.452,-3.0982,-18.597,-12.695,-75.302,-60.674,-6.1965,-54.451,-6.6386,-74.523
1027.000000000,6409.7,1198.6,1760.7,1432.1,1428.1,1180.7,2854.0,446.87,1611.3,319.09,635.33,724.37,0.0000,-3684.4,-6694.1,-313.32,-2767.4,-2660.2,-13735.,-1743.2,-1366.3,-5250.0,-2858.5,-5733.7,0.36203E+06,0.16182E+06,0.12396E+06,0.11634E+06,0.22553E+06,77716.,0.27857E+06,80500.,0.12306E+06,36733.,52792.,63591.,0.0000,-373.07,-387.20,-58.609,-352.19,-240.61,-1424.5,-1148.2,-117.22,-1030.1,-125.58,-1409.7
1028.000000000,6393.2,1292.4,1826.6,1447.9,1483.5,1293.3,3016.3,469.34,1604.1,336.05,671.64,760.75,0.0000,-3703.8,-6715.3,-315.65,-2768.7,-2672.0,-13740.,-1751.5,-1375.0,-5260.6,-2861.0,-5746.2,0.15883E+06,70993.,54382.,51040.,98942.,34095.,0.12221E+06,35316.,53990.,16115.,23161.,27898.,0.0000,-164.54,-170.21,-25.713,-154.99,-106.54,-626.20,-504.24,-51.425,-452.14,-55.146,-619.29
1029.000000000,6415.1,1367.8,1841.2,1458.6,1513.0,1285.7,3029.3,475.50,1604.7,358.36,707.70,780.69,0.0000,-3679.7,-6715.0,-313.61,-2770.7,-2654.1,-13747.,-1735.6,-1359.2,-5256.7,-2863.6,-5741.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1030.000000000,6552.6,1424.1,1785.9,1469.9,1521.4,1219.0,2962.2,475.72,1597.0,351.11,738.97,802.88,0.0000,-3674.8,-6705.9,-311.52,-2773.0,-2649.3,-13750.,-1723.2,-1352.0,-5254.7,-2868.8,-5737.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1031.000000000,6589.7,1412.2,1803.3,1470.6,1524.7,1166.6,2953.3,496.52,1604.8,332.84,785.28,781.52,0.0000,-3669.1,-6700.3,-310.04,-2772.7,-2645.1,-13752.,-1714.0,-1347.8,-5250.9,-2875.5,-5733.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1032.000000000,6659.5,1420.5,1782.1,1465.5,1556.8,1143.8,2924.5,500.13,1611.0,326.67,780.18,775.75,0.0000,-3665.3,-6693.1,-309.02,-2771.5,-2641.6,-13754.,-1707.5,-1344.5,-5246.2,-2880.1,-5730.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1033.000000000,6720.3,1379.7,1783.5,1456.9,1534.4,1171.8,3024.4,506.24,1635.8,326.69,741.76,747.83,0.0000,-3706.8,-6707.5,-312.32,-2770.1,-2665.6,-13757.,-1704.9,-1364.0,-5254.4,-2882.3,-5735.4,14152.,6325.8,4845.7,4547.9,8816.2,3038.0,10890.,3146.9,4810.8,1436.0,2063.7,2485.9,0.0000,-14.673,-15.170,-2.2911,-13.813,-9.4806,-55.846,-44.994,-4.5822,-40.323,-4.9195,-55.279
1034.000000000,6742.9,1388.9,1758.7,1455.0,1551.5,1165.7,3036.0,498.75,1611.8,334.23,705.84,755.22,0.0000,-3727.2,-6723.5,-315.61,-2769.2,-2673.0,-13759.,-1729.8,-1376.0,-5261.5,-2881.1,-5744.0,0.21129E+06,94443.,72346.,67899.,0.13162E+06,45357.,0.16258E+06,46982.,71824.,21439.,30811.,37113.,0.0000,-219.45,-226.62,-34.206,-206.42,-141.71,-833.54,-671.91,-68.412,-602.02,-73.434,-825.32
1035.000000000,6728.7,1384.9,1821.8,1449.6,1574.1,1174.8,3054.0,495.87,1617.1,341.25,690.51,766.83,0.0000,-3698.5,-6716.7,-314.24,-2768.7,-2651.5,-13760.,-1720.1,-1361.5,-5252.3,-2876.3,-5739.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1036.000000000,6750.4,1430.1,1867.3,1456.6,1660.4,1207.9,3036.2,501.31,1608.1,350.96,725.69,775.96,0.0000,-3692.8,-6710.2,-312.59,-2769.1,-2648.8,-13764.,-1712.5,-1354.8,-5249.3,-2876.0,-5737.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1037.000000000,6709.0,1389.6,1834.8,1453.0,1611.6,1185.3,2950.3,496.02,1610.8,347.63,728.46,770.23,0.0000,-3687.0,-6701.0,-311.24,-2769.9,-2645.7,-13765.,-1706.8,-1350.3,-5247.5,-2878.0,-5734.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1038.000000000,6511.0,1362.2,1803.5,1457.8,1553.5,1169.3,2982.6,495.73,1628.5,348.20,707.10,790.38,0.0000,-3681.2,-6693.9,-310.18,-2770.2,-2642.0,-13765.,-1702.7,-1347.1,-5246.1,-2878.6,-5733.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1039.000000000,6434.6,1342.5,1849.8,1488.8,1591.8,1162.4,2926.8,490.95,1617.3,339.54,692.11,778.87,0.0000,-3676.8,-6686.3,-309.37,-2770.5,-2638.6,-13764.,-1699.8,-1345.2,-5243.5,-2878.0,-5731.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1040.000000000,6287.4,1352.6,1878.1,1487.1,1597.0,1158.6,2945.8,487.87,1601.6,341.24,702.17,769.69,0.0000,-3672.2,-6680.2,-308.72,-2770.3,-2636.1,-13765.,-1697.7,-1342.9,-5242.1,-2878.2,-5729.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1041.000000000,6276.7,1361.4,1895.7,1486.3,1658.0,1164.7,2953.7,486.62,1589.5,350.68,704.29,756.28,0.0000,-3713.1,-6699.1,-312.24,-2771.1,-2661.9,-13766.,-1697.6,-1362.8,-5253.3,-2881.2,-5736.6,8892.1,3974.6,3044.6,2857.5,5539.4,1908.8,6842.2,1977.2,3022.7,902.23,1296.7,1561.9,0.0000,-9.2262,-9.5399,-1.4395,-8.6852,-5.9506,-35.092,-28.292,-2.8791,-25.347,-3.0892,-34.761
1042.000000000,6253.7,1370.2,1903.6,1482.8,1650.6,1182.9,2938.7,489.00,1598.6,349.44,695.64,749.61,0.0000,-3733.4,-6719.0,-315.63,-2772.3,-2671.0,-13767.,-1697.4,-1375.2,-5256.2,-2881.4,-5738.8,8034.1,3591.1,2750.9,2581.8,5004.9,1724.6,6181.9,1786.4,2731.0,815.18,1171.6,1411.2,0.0000,-8.3534,-8.6251,-1.3006,-7.8570,-5.3908,-31.705,-25.561,-2.6013,-22.902,-2.7910,-31.406
1043.000000000,6214.5,1374.1,1905.8,1511.4,1615.3,1187.9,2959.4,489.08,1591.1,353.55,678.93,744.09,0.0000,-3705.4,-6714.6,-314.27,-2773.2,-2649.4,-13766.,-1696.2,-1361.1,-5245.3,-2877.6,-5731.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1044.000000000,6201.0,1376.5,1907.1,1543.4,1589.4,1184.0,2980.8,485.84,1582.8,357.36,669.39,737.07,0.0000,-3696.8,-6706.6,-312.52,-2774.0,-2643.7,-13766.,-1695.2,-1354.5,-5242.0,-2874.8,-5728.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1045.000000000,6208.6,1361.4,1932.9,1555.4,1594.6,1196.6,2958.1,477.12,1594.5,359.75,672.12,745.26,0.0000,-3690.4,-6699.5,-311.10,-2775.3,-2640.9,-13766.,-1694.5,-1350.0,-5240.7,-2873.0,-5727.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1046.000000000,6300.8,1338.1,1973.4,1552.1,1593.1,1183.6,2931.7,480.64,1569.6,355.25,675.53,739.86,0.0000,-3684.7,-6692.8,-310.01,-2776.7,-2638.6,-13766.,-1694.0,-1346.5,-5239.8,-2872.3,-5726.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1047.000000000,6310.7,1315.9,1976.1,1544.9,1590.5,1179.9,2919.3,478.94,1561.3,350.31,677.22,737.67,0.0000,-3679.2,-6686.9,-309.16,-2777.9,-2636.5,-13765.,-1693.6,-1343.5,-5239.1,-2872.2,-5726.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1048.000000000,6328.1,1341.1,1959.6,1553.2,1547.9,1208.6,2938.9,484.90,1557.6,346.20,683.40,738.65,0.0000,-3719.3,-6704.9,-312.54,-2779.2,-2662.5,-13766.,-1693.9,-1363.1,-5249.8,-2874.8,-5733.6,4389.8,1962.1,1503.1,1410.7,2734.6,942.34,3377.8,976.10,1492.2,445.41,640.13,771.07,0.0000,-4.5557,-4.7114,-0.71066,-4.2886,-2.9319,-17.312,-13.959,-1.4213,-12.510,-1.5238,-17.147
1049.000000000,6307.3,1372.0,1960.6,1559.3,1543.3,1201.8,2961.7,484.97,1576.2,349.25,673.97,730.06,0.0000,-3738.6,-6725.4,-315.86,-2780.8,-2671.8,-13766.,-1695.7,-1375.6,-5253.8,-2875.4,-5736.5,15275.,6827.8,5230.3,4908.8,9515.9,3279.1,11754.,3396.6,5192.6,1549.9,2227.5,2683.1,0.0000,-15.886,-16.405,-2.4729,-14.942,-10.230,-60.240,-48.569,-4.9459,-43.529,-5.3028,-59.659
1050.000000000,6296.0,1378.2,1910.8,1550.9,1540.0,1197.6,2969.3,486.51,1576.3,352.92,671.24,711.58,0.0000,-3754.6,-6744.0,-318.58,-2782.4,-2678.7,-13767.,-1695.3,-1385.3,-5255.2,-2874.8,-5737.3,2768.1,1237.3,947.79,889.53,1724.4,594.21,2129.9,615.50,940.95,280.86,403.65,486.22,0.0000,-2.8849,-2.9750,-0.44813,-2.7106,-1.8581,-10.916,-8.8004,-0.89625,-7.8875,-0.96096,-10.810
1051.000000000,6285.7,1368.2,1907.1,1560.7,1560.5,1194.2,2939.7,489.01,1553.3,352.61,663.64,705.53,0.0000,-3768.7,-6760.1,-320.76,-2784.1,-2685.1,-13768.,-1695.3,-1392.9,-5255.9,-2874.2,-5737.5,5040.5,2253.0,1725.9,1619.8,3140.0,1082.0,3878.5,1120.8,1713.4,511.44,735.02,885.38,0.0000,-5.2643,-5.4217,-0.81601,-4.9409,-3.3909,-19.876,-16.024,-1.6320,-14.362,-1.7499,-19.682
1052.000000000,6196.2,1328.3,1739.3,1549.7,1520.6,1197.6,2907.8,492.81,1554.5,352.30,653.39,705.92,0.0000,-3735.6,-6750.9,-318.48,-2785.4,-2663.0,-13768.,-1694.6,-1375.3,-5244.1,-2871.3,-5729.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1053.000000000,6138.8,1321.8,1775.0,1520.9,1517.2,1195.2,2928.9,499.10,1545.5,344.11,649.73,711.09,0.0000,-3723.6,-6740.3,-316.12,-2785.6,-2657.2,-13768.,-1693.9,-1367.0,-5239.5,-2870.0,-5726.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1054.000000000,6126.8,1307.0,1764.4,1492.7,1518.1,1188.2,2915.9,505.69,1559.8,346.08,655.32,713.74,0.0000,-3714.4,-6729.2,-314.28,-2785.7,-2653.3,-13768.,-1693.5,-1361.4,-5237.4,-2868.8,-5725.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1055.000000000,6096.1,1301.7,1737.6,1484.2,1506.2,1175.5,2894.1,504.55,1546.3,352.13,658.21,717.06,0.0000,-3706.4,-6718.2,-312.89,-2785.4,-2649.7,-13768.,-1693.1,-1356.9,-5236.5,-2867.8,-5724.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1056.000000000,6079.3,1289.7,1698.7,1494.2,1499.8,1157.0,2879.0,503.33,1541.6,353.08,652.94,727.72,0.0000,-3699.3,-6708.7,-311.84,-2784.8,-2646.0,-13769.,-1692.8,-1353.1,-5235.8,-2866.4,-5724.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1057.000000000,6041.6,1286.7,1666.2,1513.1,1498.2,1137.6,2852.6,501.44,1557.8,354.92,645.39,728.72,0.0000,-3692.9,-6700.6,-311.02,-2784.4,-2642.9,-13769.,-1692.6,-1349.8,-5235.4,-2864.9,-5723.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1058.000000000,6030.9,1270.5,1702.9,1548.5,1515.0,1133.4,2782.7,504.47,1564.4,355.93,640.23,727.79,0.0000,-3686.9,-6693.6,-310.35,-2784.2,-2639.9,-13768.,-1692.4,-1346.6,-5235.2,-2863.7,-5722.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1059.000000000,6029.2,1228.9,1712.0,1568.0,1531.0,1123.3,2780.4,506.51,1589.8,351.14,629.98,724.81,0.0000,-3681.2,-6687.5,-309.80,-2783.9,-2637.1,-13767.,-1692.3,-1343.7,-5234.6,-2862.3,-5722.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1060.000000000,6245.2,1257.5,1728.6,1566.5,1600.9,1158.9,2785.0,493.90,1595.1,351.81,618.60,727.41,0.0000,-3720.6,-6704.7,-313.38,-2783.9,-2662.3,-13766.,-1693.1,-1363.0,-5245.7,-2863.7,-5730.1,6536.5,2921.7,2238.1,2100.5,4072.0,1403.2,5029.6,1453.4,2222.0,663.23,953.18,1148.1,0.0000,-6.7870,-7.0232,-1.0582,-6.3954,-4.3637,-25.754,-20.762,-2.1164,-18.617,-2.2685,-25.496
1061.000000000,6352.0,1282.3,1713.7,1538.6,1628.1,1187.3,2788.4,487.86,1582.9,354.51,609.27,722.23,0.0000,-3738.8,-6722.6,-316.83,-2784.0,-2670.7,-13766.,-1697.1,-1375.0,-5249.8,-2863.8,-5734.0,31216.,13953.,10688.,10031.,19446.,6701.1,24020.,6941.1,10611.,3167.3,4552.0,5483.1,0.0000,-32.474,-33.560,-5.0536,-30.576,-20.896,-122.98,-99.146,-10.107,-88.908,-10.834,-121.75
1062.000000000,6392.8,1293.2,1700.2,1537.7,1744.0,1195.1,2855.9,486.37,1558.4,357.89,593.64,723.81,0.0000,-3753.0,-6738.9,-319.61,-2784.3,-2676.8,-13767.,-1713.4,-1384.1,-5254.8,-2863.7,-5740.6,0.13132E+06,58696.,44963.,42199.,81804.,28189.,0.10104E+06,29199.,44638.,13324.,19149.,23066.,0.0000,-136.87,-141.28,-21.259,-128.74,-88.108,-517.30,-417.11,-42.518,-374.01,-45.574,-512.12
1063.000000000,6381.3,1286.3,1691.9,1558.0,1730.2,1220.5,2896.8,485.66,1567.1,355.33,593.60,705.45,0.0000,-3765.8,-6753.9,-321.81,-2784.5,-2682.2,-13770.,-1708.8,-1391.9,-5256.7,-2863.5,-5743.5,5645.7,2523.5,1933.1,1814.3,3517.0,1212.0,4344.2,1255.4,1919.2,572.84,823.28,991.68,0.0000,-5.8960,-6.0788,-0.91399,-5.5395,-3.7962,-22.240,-17.933,-1.8280,-16.080,-1.9594,-22.017
1064.000000000,6482.9,1279.5,1698.2,1534.7,1661.9,1221.7,2927.7,486.07,1557.9,359.41,587.42,708.85,0.0000,-3732.2,-6743.9,-319.50,-2784.6,-2660.0,-13771.,-1704.1,-1374.9,-5245.0,-2860.9,-5735.8,24.946,11.150,8.5416,8.0166,15.540,5.3551,19.195,5.5470,8.4800,2.5312,3.6377,4.3818,0.0000,-0.26043E-01,-0.26869E-01,-0.40386E-02,-0.24462E-01,-0.16753E-01,-0.98292E-01,-0.79243E-01,-0.80771E-02,-0.71052E-01,-0.86570E-02,-0.97303E-01
1065.000000000,6501.5,1307.9,1706.7,1518.0,1635.8,1273.6,2958.3,480.99,1552.4,357.65,603.41,704.93,0.0000,-3721.2,-6731.8,-317.11,-2784.8,-2654.9,-13774.,-1700.6,-1367.2,-5240.5,-2860.3,-5732.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1066.000000000,6469.7,1319.9,1689.0,1526.4,1604.7,1257.0,2971.9,481.50,1522.3,354.33,608.50,704.03,0.0000,-3713.0,-6721.1,-315.23,-2784.6,-2651.0,-13776.,-1698.0,-1361.9,-5238.1,-2859.8,-5729.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1067.000000000,6236.4,1292.8,1660.4,1540.8,1564.5,1241.9,2918.9,482.09,1539.4,351.64,608.57,712.01,0.0000,-3705.0,-6710.6,-313.78,-2784.8,-2647.2,-13776.,-1696.2,-1357.7,-5236.7,-2859.0,-5727.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1068.000000000,6212.3,1264.2,1691.9,1509.3,1534.1,1260.8,2850.5,480.19,1539.4,350.71,607.37,711.51,0.0000,-3698.0,-6700.9,-312.65,-2785.3,-2643.9,-13775.,-1694.9,-1354.0,-5235.0,-2858.7,-5726.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1069.000000000,6130.0,1253.4,1687.4,1498.4,1611.6,1237.3,2822.5,475.23,1518.9,346.98,608.16,721.62,0.0000,-3691.7,-6692.6,-311.74,-2785.6,-2640.8,-13773.,-1694.0,-1350.6,-5233.6,-2858.2,-5724.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1070.000000000,6046.8,1254.5,1700.8,1506.3,1620.8,1202.1,2768.6,472.51,1498.5,350.82,604.07,723.90,0.0000,-3685.4,-6685.2,-310.98,-2786.0,-2637.6,-13771.,-1693.4,-1347.4,-5232.5,-2857.3,-5723.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1071.000000000,6020.8,1221.7,1751.1,1529.5,1637.7,1202.3,2749.6,471.57,1477.7,350.56,609.35,714.52,0.0000,-3679.2,-6677.7,-310.33,-2787.1,-2634.8,-13769.,-1692.9,-1344.7,-5231.8,-2856.7,-5723.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1072.000000000,6057.8,1256.7,1761.7,1542.8,1996.2,1176.2,2776.5,475.18,1476.6,349.86,625.60,703.72,0.0000,-3673.6,-6671.1,-309.77,-2787.8,-2632.0,-13767.,-1692.5,-1342.3,-5231.0,-2856.3,-5722.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1073.000000000,6056.1,1279.0,1791.5,1545.2,1969.7,1175.3,2795.5,481.33,1463.0,351.98,636.44,707.92,0.0000,-3668.3,-6666.0,-309.27,-2788.1,-2629.4,-13766.,-1692.3,-1340.2,-5230.3,-2856.1,-5721.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1074.000000000,6029.5,1280.8,1806.8,1534.5,1916.8,1174.8,2845.6,480.41,1462.4,352.60,631.76,699.29,0.0000,-3663.1,-6661.1,-308.83,-2787.7,-2626.8,-13764.,-1692.1,-1338.4,-5229.8,-2856.0,-5720.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1075.000000000,6032.7,1240.2,1783.8,1498.7,1890.0,1209.7,2889.8,486.69,1493.9,361.32,628.34,701.76,0.0000,-3658.1,-6656.6,-308.42,-2786.7,-2624.4,-13762.,-1691.9,-1336.4,-5229.3,-2855.7,-5719.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1076.000000000,6073.9,1217.4,1767.1,1481.0,1746.9,1231.0,2849.6,493.22,1466.7,357.91,624.98,714.06,0.0000,-3653.2,-6653.7,-308.03,-2785.7,-2621.9,-13760.,-1691.8,-1334.5,-5229.2,-2855.7,-5719.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1077.000000000,6043.8,1206.0,1738.7,1477.3,1632.4,1232.0,2792.6,491.28,1471.9,356.21,626.67,713.27,0.0000,-3693.1,-6676.1,-311.70,-2784.9,-2647.5,-13759.,-1712.3,-1354.1,-5244.5,-2857.9,-5732.3,0.15405E+06,68857.,52746.,49504.,95966.,33069.,0.11854E+06,34254.,52366.,15631.,22464.,27059.,0.0000,-159.36,-165.18,-24.939,-150.49,-102.25,-607.05,-489.16,-49.878,-438.68,-53.440,-600.43
1078.000000000,6004.2,1209.1,1717.0,1468.7,1738.3,1192.9,2756.6,496.35,1446.2,353.60,621.08,727.11,0.0000,-3667.3,-6676.1,-311.12,-2784.1,-2628.4,-13757.,-1707.1,-1344.6,-5237.6,-2855.8,-5729.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1079.000000000,5939.8,1218.7,1717.6,1477.7,1754.5,1197.1,2770.0,501.27,1471.1,341.93,617.29,725.91,0.0000,-3659.8,-6669.6,-310.02,-2783.2,-2624.3,-13755.,-1702.7,-1340.3,-5234.3,-2854.5,-5727.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1080.000000000,5969.3,1218.5,1735.2,1489.1,1739.1,1205.7,2828.1,505.46,1472.5,342.57,615.13,722.39,0.0000,-3655.0,-6662.9,-309.04,-2782.8,-2622.6,-13754.,-1699.4,-1337.5,-5231.8,-2853.8,-5725.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1081.000000000,5959.1,1229.8,1757.7,1489.9,1732.2,1205.6,2850.4,509.83,1452.4,345.96,631.12,714.37,0.0000,-3651.4,-6657.9,-308.26,-2782.2,-2620.7,-13754.,-1697.0,-1335.1,-5229.8,-2853.2,-5723.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1082.000000000,5799.6,1257.4,1750.7,1470.5,1713.2,1169.8,2803.4,508.50,1425.9,348.32,614.75,720.37,0.0000,-3647.1,-6653.4,-307.60,-2781.3,-2617.8,-13754.,-1695.3,-1332.8,-5228.8,-2852.2,-5721.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1083.000000000,5811.6,1250.8,1718.8,1483.9,1745.7,1155.9,2761.3,489.77,1443.9,353.57,601.60,728.13,0.0000,-3642.2,-6648.2,-307.03,-2780.6,-2615.1,-13753.,-1694.1,-1330.8,-5227.5,-2851.4,-5720.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1084.000000000,5973.4,1233.9,1709.3,1475.1,1777.2,1179.0,2744.3,485.06,1466.6,347.56,602.37,731.32,0.0000,-3637.8,-6643.9,-306.53,-2780.1,-2612.5,-13751.,-1693.3,-1329.0,-5226.3,-2851.2,-5718.9,19.637,8.7774,6.7237,6.3105,12.233,4.2155,15.110,4.3665,6.6753,1.9925,2.8636,3.4493,0.0000,-0.20218E-01,-0.21012E-01,-0.31791E-02,-0.19145E-01,-0.12977E-01,-0.77411E-01,-0.62354E-01,-0.63581E-02,-0.55920E-01,-0.68099E-02,-0.76534E-01
1085.000000000,5825.9,1240.3,1743.5,1465.4,1769.5,1184.0,2727.4,489.33,1479.6,347.99,592.78,737.23,0.0000,-3633.4,-6640.0,-306.08,-2779.2,-2610.1,-13750.,-1692.7,-1327.4,-5225.4,-2850.4,-5718.1,5.4414,2.4322,1.8631,1.7486,3.3898,1.1681,4.1870,1.2099,1.8497,0.55211,0.79348,0.95579,0.0000,-0.55979E-02,-0.58200E-02,-0.88092E-03,-0.53035E-02,-0.35932E-02,-0.21448E-01,-0.17277E-01,-0.17618E-02,-0.15495E-01,-0.18869E-02,-0.21206E-01
1086.000000000,5757.3,1264.5,1767.3,1478.2,1740.4,1181.2,2784.3,497.44,1499.1,345.98,595.34,730.23,0.0000,-3629.3,-6637.1,-305.69,-2778.3,-2607.8,-13750.,-1692.2,-1326.0,-5224.5,-2850.2,-5717.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1087.000000000,5824.8,1262.8,1743.1,1471.4,1777.3,1176.7,2765.2,491.29,1503.7,345.40,602.60,729.97,0.0000,-3625.5,-6634.4,-305.32,-2777.1,-2605.5,-13749.,-1691.9,-1324.6,-5223.6,-2849.9,-5716.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1088.000000000,5774.5,1258.4,1757.0,1448.3,1765.1,1153.1,2736.4,495.70,1478.7,345.69,599.09,738.36,0.0000,-3621.9,-6632.4,-304.96,-2775.9,-2603.3,-13748.,-1691.6,-1323.4,-5222.7,-2849.7,-5716.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1089.000000000,5995.9,1250.4,1764.6,1454.3,1741.2,1156.9,2706.7,492.51,1457.5,345.53,601.44,731.61,0.0000,-3618.2,-6630.2,-304.61,-2774.7,-2600.9,-13748.,-1691.4,-1322.2,-5222.0,-2849.3,-5716.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1090.000000000,5808.1,1251.3,1754.6,1460.6,1759.0,1149.9,2719.5,493.45,1486.1,344.48,603.98,729.42,0.0000,-3614.0,-6627.7,-304.26,-2773.7,-2598.4,-13746.,-1691.3,-1321.1,-5221.3,-2848.7,-5715.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1091.000000000,5726.7,1281.1,1750.8,1458.3,1778.9,1165.3,2740.1,498.99,1488.0,341.92,599.91,737.25,0.0000,-3654.0,-6647.7,-307.94,-2772.9,-2624.0,-13746.,-1708.7,-1340.4,-5235.8,-2850.7,-5727.8,0.13056E+06,58360.,44705.,41957.,81336.,28028.,0.10047E+06,29032.,44383.,13248.,19039.,22934.,0.0000,-133.99,-139.39,-21.137,-127.10,-85.997,-514.18,-414.46,-42.274,-371.73,-45.260,-508.50
1092.000000000,5689.7,1265.1,1732.6,1463.8,1729.3,1193.7,2733.4,498.61,1491.4,341.15,600.84,731.98,0.0000,-3673.0,-6669.4,-311.45,-2772.5,-2633.0,-13746.,-1707.9,-1353.6,-5241.2,-2851.4,-5733.6,26778.,11969.,9168.7,8605.1,16681.,5748.3,20605.,5954.2,9102.6,2717.0,3904.8,4703.6,0.0000,-27.537,-28.604,-4.3351,-26.099,-17.655,-105.44,-85.003,-8.6701,-76.238,-9.2824,-104.28
1093.000000000,5745.1,1261.2,1705.9,1462.7,1727.5,1168.8,2739.6,499.93,1479.3,338.85,602.14,729.36,0.0000,-3643.9,-6666.4,-310.20,-2771.8,-2611.7,-13744.,-1703.3,-1341.8,-5230.9,-2849.4,-5727.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1094.000000000,5761.7,1266.8,1713.3,1471.9,1707.6,1155.8,2750.2,499.65,1475.4,337.83,597.91,734.93,0.0000,-3634.7,-6659.6,-308.56,-2770.8,-2606.7,-13743.,-1699.7,-1336.6,-5226.7,-2848.6,-5724.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1095.000000000,5781.1,1263.3,1723.8,1473.4,1710.5,1159.3,2768.0,503.05,1451.1,336.25,600.48,735.99,0.0000,-3628.7,-6653.1,-307.23,-2770.0,-2604.0,-13743.,-1697.0,-1333.2,-5224.3,-2848.0,-5722.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1096.000000000,5796.9,1257.1,1722.8,1463.6,1709.2,1156.9,2777.8,500.32,1459.3,334.72,601.17,733.62,0.0000,-3624.4,-6647.6,-306.22,-2769.2,-2601.8,-13742.,-1695.1,-1330.6,-5222.6,-2847.4,-5720.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1097.000000000,5913.8,1256.9,1735.4,1484.1,1696.2,1183.0,2778.5,500.49,1466.1,335.10,600.60,734.13,0.0000,-3664.6,-6666.6,-309.47,-2768.4,-2627.4,-13743.,-1694.1,-1349.6,-5232.8,-2849.3,-5727.5,1700.1,759.90,582.10,546.32,1059.1,364.95,1308.1,378.02,577.90,172.50,247.91,298.62,0.0000,-1.7485,-1.8160,-0.27523,-1.6564,-1.1198,-6.6936,-5.3966,-0.55045,-4.8404,-0.58930,-6.6207
1098.000000000,5930.2,1251.3,1732.5,1497.5,1690.7,1204.0,2804.2,499.11,1476.1,336.15,596.26,727.97,0.0000,-3683.4,-6687.5,-312.70,-2767.7,-2636.0,-13743.,-1696.4,-1362.1,-5236.3,-2849.7,-5730.2,23738.,10611.,8128.0,7628.4,14788.,5095.8,18266.,5278.4,8069.4,2408.6,3461.6,4169.7,0.0000,-24.463,-25.371,-3.8430,-23.153,-15.653,-93.453,-75.354,-7.6860,-67.587,-8.2284,-92.442
1099.000000000,5929.1,1230.9,1724.1,1501.3,1677.0,1190.0,2804.0,499.25,1467.5,337.04,596.99,730.06,0.0000,-3653.7,-6683.0,-311.26,-2766.9,-2614.4,-13742.,-1694.9,-1349.1,-5225.7,-2847.1,-5723.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1100.000000000,5909.7,1230.3,1707.7,1510.3,1606.8,1176.0,2808.5,501.43,1459.9,335.49,595.35,729.74,0.0000,-3644.1,-6674.9,-309.47,-2766.3,-2608.8,-13741.,-1693.7,-1343.1,-5222.1,-2846.1,-5720.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1101.000000000,5906.1,1226.9,1698.1,1521.4,1574.6,1170.8,2795.4,497.89,1452.0,334.49,592.66,730.61,0.0000,-3637.4,-6666.8,-308.00,-2765.6,-2605.1,-13740.,-1692.8,-1339.1,-5220.4,-2845.3,-5718.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1102.000000000,5797.0,1235.7,1698.9,1519.2,1550.2,1174.1,2791.6,498.26,1455.9,333.29,592.75,730.69,0.0000,-3631.3,-6659.2,-306.86,-2764.9,-2601.9,-13739.,-1692.1,-1335.7,-5219.3,-2844.4,-5717.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1103.000000000,5722.5,1230.3,1707.1,1515.5,1540.1,1177.6,2781.4,498.53,1457.2,332.59,592.55,729.55,0.0000,-3625.8,-6652.7,-305.96,-2764.2,-2599.1,-13738.,-1691.6,-1332.7,-5218.2,-2843.7,-5717.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1104.000000000,5713.5,1219.8,1722.2,1510.5,1526.7,1174.9,2782.7,500.62,1467.7,331.71,588.19,724.98,0.0000,-3620.8,-6646.6,-305.23,-2763.5,-2596.5,-13736.,-1691.2,-1330.1,-5217.2,-2843.1,-5716.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1105.000000000,5722.0,1225.1,1720.7,1511.3,1527.3,1168.9,2781.1,505.01,1470.4,332.54,583.68,727.67,0.0000,-3616.0,-6641.4,-304.61,-2762.7,-2594.0,-13735.,-1690.9,-1327.7,-5216.7,-2842.6,-5716.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1106.000000000,5736.5,1211.8,1712.9,1513.9,1554.8,1166.2,2745.8,506.71,1479.5,332.61,583.35,725.77,0.0000,-3611.5,-6637.3,-304.09,-2761.9,-2591.6,-13735.,-1690.7,-1325.7,-5216.2,-2842.0,-5715.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1107.000000000,5762.9,1209.1,1700.1,1511.4,1556.8,1161.8,2727.9,504.86,1478.1,334.26,586.97,721.51,0.0000,-3607.1,-6633.7,-303.63,-2761.0,-2589.1,-13734.,-1690.5,-1323.9,-5215.7,-2841.6,-5715.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1108.000000000,5721.9,1219.0,1708.3,1518.7,1556.3,1159.5,2716.4,502.61,1472.4,331.48,584.96,715.74,0.0000,-3602.9,-6630.1,-303.21,-2760.2,-2586.7,-13732.,-1690.3,-1322.3,-5215.2,-2840.9,-5715.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1109.000000000,5636.3,1217.4,1724.7,1530.4,1563.9,1176.1,2711.7,502.22,1466.3,331.04,584.08,712.40,0.0000,-3599.0,-6626.5,-302.83,-2759.4,-2584.5,-13731.,-1690.2,-1320.7,-5214.8,-2840.2,-5714.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1110.000000000,5635.0,1219.7,1719.3,1535.0,1552.1,1172.0,2712.0,503.31,1476.4,329.88,584.54,708.73,0.0000,-3595.3,-6622.2,-302.46,-2758.7,-2582.4,-13730.,-1690.1,-1319.2,-5214.3,-2839.5,-5714.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1111.000000000,5646.4,1205.5,1712.6,1538.8,1539.6,1173.5,2700.5,505.53,1477.3,330.20,582.59,705.66,0.0000,-3591.8,-6618.2,-302.10,-2758.1,-2580.4,-13729.,-1690.0,-1317.8,-5214.0,-2839.0,-5714.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1112.000000000,5515.5,1199.4,1704.6,1552.1,1532.5,1182.1,2684.5,504.87,1486.4,329.78,580.34,706.24,0.0000,-3588.3,-6614.8,-301.76,-2757.5,-2578.4,-13728.,-1689.9,-1316.5,-5213.6,-2838.5,-5714.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1113.000000000,5458.0,1203.0,1700.4,1561.0,1527.3,1197.9,2682.9,505.56,1486.7,329.14,575.96,706.39,0.0000,-3585.1,-6611.8,-301.43,-2756.9,-2576.4,-13727.,-1689.8,-1315.4,-5213.1,-2837.8,-5714.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1114.000000000,5472.0,1194.9,1695.2,1561.8,1517.8,1192.6,2673.9,502.32,1485.1,327.37,576.16,702.52,0.0000,-3582.2,-6609.0,-301.10,-2756.2,-2574.5,-13726.,-1689.7,-1314.2,-5212.6,-2837.1,-5713.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1115.000000000,5464.0,1179.0,1692.1,1576.7,1503.9,1190.6,2661.1,504.57,1485.2,327.91,573.23,697.81,0.0000,-3579.1,-6606.8,-300.78,-2755.5,-2572.5,-13725.,-1689.6,-1313.2,-5212.1,-2836.4,-5713.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1116.000000000,5269.3,1177.4,1674.4,1569.7,1523.6,1193.5,2639.0,506.03,1497.2,326.14,570.68,695.08,0.0000,-3575.8,-6604.7,-300.47,-2754.7,-2570.6,-13724.,-1689.5,-1312.2,-5211.6,-2835.6,-5713.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1117.000000000,5205.9,1177.9,1665.7,1565.8,1589.8,1204.6,2647.7,508.36,1492.1,326.68,569.05,693.56,0.0000,-3572.7,-6602.4,-300.16,-2753.9,-2568.8,-13722.,-1689.5,-1311.2,-5211.1,-2834.9,-5713.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1118.000000000,5285.0,1169.2,1672.3,1567.2,1611.5,1209.4,2657.0,508.33,1476.0,325.16,563.16,689.16,0.0000,-3569.7,-6600.2,-299.85,-2753.3,-2567.0,-13721.,-1689.4,-1310.3,-5210.6,-2834.1,-5712.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1119.000000000,5336.5,1162.9,1681.4,1574.2,1610.5,1201.3,2669.6,504.70,1488.5,324.99,558.32,680.58,0.0000,-3566.7,-6598.0,-299.54,-2752.8,-2565.5,-13720.,-1689.3,-1309.6,-5210.2,-2833.4,-5712.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1120.000000000,5335.7,1156.1,1683.6,1584.1,1597.7,1190.7,2651.4,500.31,1476.1,327.37,558.80,682.53,0.0000,-3563.6,-6596.0,-299.24,-2752.3,-2563.9,-13718.,-1689.2,-1308.8,-5209.8,-2833.0,-5712.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1121.000000000,5339.5,1156.6,1681.9,1594.4,1605.5,1196.3,2632.5,500.25,1466.8,326.01,560.59,685.95,0.0000,-3560.6,-6594.0,-298.94,-2751.7,-2562.3,-13717.,-1689.1,-1308.1,-5209.4,-2832.6,-5711.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1122.000000000,5358.2,1153.3,1700.4,1595.2,1601.8,1210.6,2603.7,498.59,1490.0,323.37,565.58,688.06,0.0000,-3601.5,-6615.2,-302.65,-2751.2,-2588.5,-13717.,-1699.8,-1326.4,-5222.7,-2834.7,-5722.4,79640.,35597.,27269.,25592.,49612.,17096.,61280.,17708.,27072.,8080.6,11613.,13989.,0.0000,-80.947,-84.427,-12.893,-77.107,-51.580,-312.70,-252.40,-25.786,-226.56,-27.551,-309.32
1123.000000000,5109.3,1149.8,1693.6,1589.4,1627.5,1211.4,2600.0,499.10,1493.4,323.42,564.75,689.08,0.0000,-3577.1,-6614.8,-302.17,-2750.7,-2570.1,-13715.,-1697.0,-1319.0,-5215.4,-2832.6,-5718.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1124.000000000,5237.3,1158.8,1688.9,1590.1,1618.6,1218.4,2599.1,499.15,1493.3,324.79,565.07,686.82,0.0000,-3570.4,-6610.8,-301.16,-2750.1,-2566.2,-13713.,-1694.8,-1315.6,-5212.8,-2831.6,-5716.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1125.000000000,5236.4,1158.2,1687.1,1586.5,1613.4,1214.4,2597.2,499.62,1492.1,326.98,565.24,688.10,0.0000,-3566.0,-6606.3,-300.25,-2749.4,-2563.8,-13712.,-1693.0,-1313.4,-5211.1,-2830.6,-5715.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1126.000000000,5239.8,1165.1,1687.3,1585.8,1615.6,1214.7,2563.0,497.97,1486.9,327.40,564.06,691.05,0.0000,-3562.1,-6602.3,-299.52,-2748.6,-2561.8,-13711.,-1691.7,-1311.7,-5209.7,-2829.8,-5713.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1127.000000000,5227.2,1172.6,1680.0,1594.6,1624.9,1205.3,2565.3,496.53,1471.3,327.41,562.78,689.67,0.0000,-3558.6,-6598.8,-298.92,-2747.8,-2559.9,-13710.,-1690.8,-1310.2,-5208.6,-2829.0,-5712.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1128.000000000,5248.7,1172.1,1676.7,1597.5,1635.9,1204.5,2554.1,493.73,1465.0,326.66,558.46,689.17,0.0000,-3555.3,-6595.7,-298.41,-2746.9,-2558.2,-13709.,-1690.1,-1308.9,-5207.7,-2828.3,-5711.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1129.000000000,5378.4,1189.1,1692.9,1591.9,1661.8,1208.9,2537.6,494.96,1465.8,324.47,547.59,687.28,0.0000,-3552.2,-6593.1,-297.98,-2746.1,-2556.5,-13708.,-1689.6,-1307.8,-5206.9,-2827.6,-5710.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1130.000000000,5372.6,1180.8,1711.2,1592.0,1671.0,1222.4,2504.5,495.33,1478.3,325.71,544.80,686.54,0.0000,-3549.3,-6590.5,-297.60,-2745.3,-2554.9,-13706.,-1689.3,-1306.7,-5206.4,-2826.8,-5710.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1131.000000000,5307.5,1162.0,1713.6,1588.1,1666.3,1228.8,2494.3,493.62,1494.9,326.66,542.18,686.93,0.0000,-3546.5,-6587.9,-297.21,-2744.6,-2553.3,-13704.,-1689.0,-1305.6,-5205.8,-2825.7,-5709.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1132.000000000,5274.2,1159.6,1724.6,1597.0,1669.2,1229.9,2511.7,494.22,1493.8,325.50,538.64,683.12,0.0000,-3543.8,-6585.6,-296.84,-2743.8,-2551.7,-13703.,-1688.8,-1304.5,-5205.3,-2824.7,-5708.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1133.000000000,5308.3,1173.7,1727.4,1575.6,1767.5,1222.7,2521.8,493.66,1496.4,324.41,540.17,681.50,0.0000,-3541.0,-6583.3,-296.48,-2743.2,-2550.1,-13702.,-1688.6,-1303.5,-5204.7,-2823.8,-5707.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1134.000000000,5359.2,1183.8,1717.8,1585.5,1833.0,1221.3,2537.5,493.33,1492.6,319.42,541.76,679.76,0.0000,-3538.3,-6581.0,-296.15,-2742.5,-2548.6,-13700.,-1688.5,-1302.5,-5204.1,-2823.1,-5707.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1135.000000000,5339.7,1189.0,1710.3,1575.2,1846.2,1226.4,2532.9,492.60,1496.2,317.81,538.86,679.83,0.0000,-3535.6,-6578.6,-295.82,-2741.9,-2547.1,-13700.,-1688.4,-1301.5,-5203.7,-2822.3,-5706.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1136.000000000,5334.2,1187.5,1710.0,1575.3,1853.5,1223.0,2532.2,492.87,1492.2,319.89,544.16,672.55,0.0000,-3533.0,-6576.5,-295.50,-2741.5,-2545.6,-13699.,-1688.2,-1300.4,-5203.2,-2821.6,-5705.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1137.000000000,5340.3,1191.8,1719.9,1574.3,1831.1,1219.0,2544.2,494.54,1493.0,320.52,545.34,668.28,0.0000,-3530.4,-6574.8,-295.19,-2741.0,-2544.2,-13698.,-1688.1,-1299.3,-5202.8,-2821.1,-5705.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1138.000000000,5335.2,1189.7,1729.4,1576.7,1863.2,1229.9,2537.8,495.50,1503.3,319.33,546.42,667.25,0.0000,-3527.8,-6573.5,-294.89,-2740.6,-2542.8,-13697.,-1688.0,-1298.4,-5202.3,-2820.5,-5704.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1139.000000000,5332.2,1190.8,1736.0,1574.3,1875.3,1232.5,2512.3,493.03,1504.3,317.68,546.04,667.28,0.0000,-3525.1,-6572.1,-294.60,-2740.1,-2541.4,-13696.,-1687.9,-1297.6,-5202.0,-2820.0,-5704.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1140.000000000,5341.5,1202.5,1724.2,1570.2,1871.5,1240.7,2514.5,491.40,1503.6,317.54,544.99,666.39,0.0000,-3522.5,-6570.5,-294.31,-2739.8,-2539.9,-13695.,-1687.8,-1296.8,-5201.5,-2819.5,-5703.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1141.000000000,5357.2,1199.4,1697.8,1561.6,1907.3,1240.6,2500.0,486.20,1516.6,318.57,546.06,665.06,0.0000,-3520.1,-6568.8,-294.03,-2739.3,-2538.5,-13694.,-1687.7,-1296.0,-5201.2,-2818.9,-5703.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1142.000000000,5364.0,1202.7,1708.5,1564.5,1969.1,1234.9,2484.1,484.95,1517.2,316.87,548.69,672.01,0.0000,-3517.8,-6567.0,-293.75,-2738.9,-2536.9,-13693.,-1687.7,-1295.3,-5200.7,-2818.3,-5702.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1143.000000000,5368.9,1207.2,1715.5,1563.6,1967.3,1229.5,2491.8,481.71,1517.9,317.53,552.16,679.34,0.0000,-3515.4,-6565.4,-293.47,-2738.2,-2535.3,-13691.,-1687.6,-1294.6,-5200.2,-2817.7,-5702.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1144.000000000,5382.2,1207.6,1717.2,1551.2,1976.2,1227.3,2490.2,481.07,1498.0,320.14,551.07,681.01,0.0000,-3512.9,-6563.8,-293.20,-2737.5,-2533.8,-13690.,-1687.5,-1294.0,-5199.8,-2817.1,-5702.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1145.000000000,5390.7,1222.1,1713.4,1549.8,1986.9,1226.2,2473.2,481.06,1490.3,321.03,550.88,685.22,0.0000,-3510.5,-6562.1,-292.92,-2736.9,-2532.3,-13689.,-1687.4,-1293.4,-5199.3,-2816.6,-5701.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1146.000000000,5401.4,1224.6,1708.8,1551.7,1986.7,1233.9,2460.1,483.19,1500.0,322.33,558.85,685.49,0.0000,-3508.1,-6560.4,-292.66,-2736.3,-2530.9,-13688.,-1687.3,-1292.8,-5198.8,-2816.1,-5701.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1147.000000000,5400.9,1227.7,1702.3,1553.8,1986.2,1234.6,2465.3,483.72,1506.1,323.97,559.63,686.01,0.0000,-3505.6,-6558.8,-292.40,-2735.7,-2529.5,-13686.,-1687.2,-1292.3,-5198.4,-2815.6,-5700.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1148.000000000,5388.0,1235.4,1704.9,1545.7,1989.2,1248.3,2463.5,480.79,1507.4,323.58,558.78,682.32,0.0000,-3546.3,-6579.9,-296.14,-2735.2,-2556.0,-13686.,-1691.2,-1309.4,-5210.3,-2817.8,-5709.5,30408.,13592.,10412.,9771.6,18943.,6527.5,23398.,6761.3,10336.,3085.3,4434.1,5341.1,0.0000,-30.613,-32.002,-4.9227,-29.293,-19.403,-119.13,-96.223,-9.8454,-86.441,-10.503,-117.81
1149.000000000,5427.0,1247.5,1708.9,1542.9,1994.7,1257.2,2490.8,483.05,1503.6,321.23,556.71,682.45,0.0000,-3566.1,-6603.0,-299.73,-2734.6,-2565.8,-13686.,-1701.5,-1322.0,-5216.3,-2818.5,-5715.4,84188.,37630.,28826.,27054.,52445.,18072.,64780.,18720.,28618.,8542.1,12277.,14788.,0.0000,-84.912,-88.662,-13.629,-81.169,-53.792,-329.82,-266.42,-27.259,-239.32,-29.080,-326.16
1150.000000000,5469.3,1248.9,1696.0,1531.7,1880.6,1247.6,2497.2,486.06,1501.3,320.47,557.36,681.10,0.0000,-3538.7,-6601.2,-298.60,-2734.0,-2545.4,-13684.,-1697.7,-1312.1,-5207.1,-2816.4,-5709.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1151.000000000,5611.7,1227.4,1699.0,1521.6,1880.6,1241.4,2502.8,485.30,1491.7,320.81,557.08,675.34,0.0000,-3531.1,-6595.4,-297.06,-2733.3,-2540.9,-13682.,-1694.7,-1307.4,-5203.8,-2815.4,-5707.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1152.000000000,5622.4,1223.2,1721.2,1520.6,1860.8,1237.2,2493.8,485.62,1484.6,323.24,554.22,673.83,0.0000,-3526.1,-6589.4,-295.79,-2732.4,-2538.3,-13681.,-1692.3,-1304.3,-5202.0,-2814.7,-5705.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1153.000000000,5768.9,1222.1,1732.9,1515.8,1900.4,1234.9,2494.9,483.54,1478.7,324.49,557.99,676.58,0.0000,-3522.0,-6584.1,-294.82,-2731.4,-2536.1,-13680.,-1690.6,-1301.8,-5200.7,-2814.2,-5703.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1154.000000000,5764.6,1228.4,1737.7,1500.1,1906.5,1239.4,2481.1,483.88,1466.5,324.26,555.82,680.14,0.0000,-3518.2,-6579.4,-294.07,-2730.6,-2534.4,-13679.,-1689.4,-1299.7,-5199.5,-2813.5,-5702.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1155.000000000,5664.3,1232.1,1741.0,1488.5,1885.2,1243.1,2481.8,483.97,1474.3,326.08,559.03,684.99,0.0000,-3515.0,-6575.4,-293.49,-2729.9,-2533.3,-13678.,-1688.6,-1297.9,-5198.5,-2813.2,-5701.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1156.000000000,5677.4,1225.0,1730.6,1495.5,1881.7,1236.1,2471.9,480.76,1480.4,323.88,563.21,686.13,0.0000,-3512.3,-6572.0,-293.02,-2729.0,-2531.6,-13677.,-1687.9,-1296.4,-5197.7,-2812.6,-5700.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1157.000000000,5680.4,1210.7,1740.5,1505.1,1892.6,1233.2,2477.6,480.88,1489.2,324.26,561.52,689.40,0.0000,-3509.3,-6569.3,-292.62,-2728.1,-2529.9,-13676.,-1687.5,-1294.9,-5197.1,-2811.9,-5699.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1158.000000000,5706.8,1211.3,1750.0,1505.4,1843.2,1234.6,2496.5,480.62,1485.8,325.34,563.36,691.36,0.0000,-3506.5,-6566.4,-292.27,-2727.2,-2528.3,-13676.,-1687.1,-1293.6,-5196.6,-2811.4,-5699.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1159.000000000,5784.7,1219.8,1762.4,1483.7,1768.6,1220.9,2511.5,480.36,1494.2,324.63,561.36,688.97,0.0000,-3503.8,-6563.8,-291.95,-2726.3,-2526.8,-13675.,-1686.9,-1292.5,-5196.1,-2810.8,-5698.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1160.000000000,5823.3,1231.2,1763.9,1483.7,1775.5,1213.5,2520.2,480.21,1500.7,324.68,553.74,686.37,0.0000,-3501.2,-6561.2,-291.65,-2725.5,-2525.2,-13674.,-1686.7,-1291.4,-5195.5,-2810.3,-5698.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1161.000000000,5813.9,1249.1,1755.9,1480.4,1779.9,1201.4,2521.1,478.12,1499.9,324.99,546.65,685.41,0.0000,-3498.7,-6559.0,-291.37,-2724.7,-2523.7,-13674.,-1686.5,-1290.3,-5194.9,-2809.8,-5697.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1162.000000000,5819.2,1256.2,1729.3,1472.0,1769.2,1200.7,2520.5,478.97,1506.1,324.97,546.87,686.46,0.0000,-3496.3,-6556.1,-291.11,-2723.8,-2522.3,-13673.,-1686.3,-1289.4,-5194.5,-2809.3,-5697.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1163.000000000,5818.0,1258.0,1716.0,1466.5,1763.8,1213.5,2520.7,484.73,1514.4,325.87,549.71,684.96,0.0000,-3537.3,-6576.5,-294.85,-2722.9,-2548.7,-13674.,-1705.0,-1306.3,-5209.5,-2811.4,-5709.6,0.14044E+06,62772.,48085.,45129.,87485.,30147.,0.10806E+06,31227.,47738.,14249.,20479.,24668.,0.0000,-141.18,-147.54,-22.735,-135.18,-89.136,-549.92,-444.26,-45.470,-399.15,-48.480,-543.70
1164.000000000,5822.7,1241.9,1707.7,1465.5,1748.0,1216.3,2536.7,490.48,1517.1,325.52,551.24,686.13,0.0000,-3557.4,-6599.1,-298.44,-2722.2,-2558.4,-13673.,-1712.2,-1318.6,-5217.3,-2812.4,-5717.6,89138.,39843.,30521.,28645.,55529.,19135.,68588.,19820.,30301.,9044.4,12998.,15657.,0.0000,-89.780,-93.706,-14.431,-85.868,-56.655,-349.02,-282.02,-28.861,-253.35,-30.773,-345.10
1165.000000000,5833.3,1252.8,1713.0,1474.7,1739.1,1216.4,2557.5,492.50,1519.4,326.66,550.63,679.37,0.0000,-3574.0,-6619.6,-301.32,-2721.5,-2565.8,-13674.,-1723.1,-1328.7,-5223.4,-2812.9,-5725.0,0.13299E+06,59444.,45536.,42737.,82847.,28549.,0.10233E+06,29571.,45208.,13494.,19393.,23360.,0.0000,-134.22,-139.93,-21.530,-128.22,-84.616,-520.76,-420.87,-43.060,-378.01,-45.913,-514.92
1166.000000000,5842.3,1314.8,1742.4,1486.6,1769.6,1263.0,2656.4,502.45,1534.9,337.12,563.34,701.64,0.0000,-3591.9,-6639.1,-303.66,-2722.3,-2576.2,-13676.,-1730.9,-1337.6,-5229.1,-2814.4,-5731.8,0.13192E+06,58967.,45170.,42394.,82182.,28319.,0.10151E+06,29334.,44844.,13386.,19237.,23172.,0.0000,-133.63,-139.04,-21.357,-127.49,-84.402,-517.20,-417.78,-42.714,-375.10,-45.571,-511.25
1167.000000000,5844.9,1368.1,1790.5,1485.6,1776.2,1286.0,2723.3,502.97,1551.8,354.82,596.35,729.81,0.0000,-3611.5,-6661.5,-305.63,-2723.5,-2586.5,-13682.,-1729.6,-1345.6,-5235.6,-2817.6,-5736.0,80687.,36065.,27627.,25929.,50264.,17321.,62086.,17941.,27428.,8186.9,11766.,14173.,0.0000,-82.094,-85.178,-13.062,-78.182,-51.941,-316.75,-255.73,-26.125,-229.53,-27.896,-313.02
1168.000000000,5836.8,1408.3,1775.0,1481.1,1742.2,1249.4,2675.2,498.50,1546.2,363.85,616.22,733.12,0.0000,-3585.7,-6655.4,-303.31,-2725.9,-2565.6,-13685.,-1717.6,-1330.6,-5227.2,-2820.0,-5728.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1169.000000000,5703.0,1410.2,1731.9,1460.2,1683.7,1229.0,2662.7,503.42,1561.3,355.31,627.31,748.05,0.0000,-3578.6,-6645.5,-301.04,-2726.7,-2560.6,-13687.,-1708.5,-1323.5,-5222.8,-2823.4,-5723.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1170.000000000,5723.5,1375.9,1754.6,1451.9,1680.8,1205.4,2624.3,513.62,1572.9,350.63,645.80,729.37,0.0000,-3572.6,-6636.5,-299.39,-2726.2,-2556.6,-13688.,-1702.0,-1319.0,-5219.7,-2826.6,-5718.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1171.000000000,5732.4,1403.8,1744.9,1454.7,1702.5,1186.0,2607.4,513.50,1573.8,342.54,662.47,727.01,0.0000,-3567.3,-6629.5,-298.25,-2725.0,-2553.2,-13688.,-1697.5,-1315.7,-5216.2,-2830.6,-5715.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1172.000000000,5715.7,1423.4,1740.1,1476.5,1738.1,1192.8,2622.5,511.30,1597.0,341.22,640.37,717.87,0.0000,-3607.7,-6644.4,-301.44,-2723.4,-2577.9,-13689.,-1694.7,-1333.5,-5224.5,-2834.5,-5721.0,2414.7,1079.3,826.80,775.98,1504.3,518.36,1858.1,536.93,820.84,245.01,352.12,424.15,0.0000,-2.4564,-2.5492,-0.39092,-2.3388,-1.5503,-9.4772,-7.6610,-0.78185,-6.8737,-0.83527,-9.3805
1173.000000000,5720.9,1429.2,1723.6,1473.5,1730.8,1181.6,2688.2,513.89,1610.0,339.36,629.31,706.22,0.0000,-3583.4,-6637.0,-300.64,-2722.0,-2558.0,-13690.,-1692.4,-1323.4,-5213.6,-2832.2,-5713.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1174.000000000,5731.1,1447.0,1543.2,1476.4,1792.9,1198.4,2692.1,510.07,1608.2,348.36,607.31,696.30,0.0000,-3620.7,-6650.2,-303.47,-2720.5,-2580.4,-13692.,-1699.5,-1339.4,-5223.6,-2832.3,-5721.1,64894.,29006.,22220.,20854.,40426.,13931.,49933.,14430.,22059.,6584.4,9463.0,11399.,0.0000,-66.086,-68.534,-10.506,-62.859,-41.593,-254.56,-205.88,-21.011,-184.72,-22.442,-252.06
1175.000000000,5722.5,1440.0,1572.0,1468.5,1789.7,1188.9,2670.2,502.65,1600.6,352.86,593.21,698.94,0.0000,-3594.5,-6644.1,-302.28,-2719.3,-2559.7,-13693.,-1696.2,-1328.0,-5214.6,-2828.6,-5715.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1176.000000000,5680.9,1424.2,1576.1,1461.2,1840.9,1184.6,2633.4,497.35,1594.5,352.84,577.16,690.78,0.0000,-3586.2,-6634.2,-300.77,-2718.4,-2554.2,-13693.,-1693.6,-1322.1,-5211.0,-2826.0,-5713.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1177.000000000,5695.3,1400.1,1549.9,1456.3,1839.6,1185.6,2629.5,496.97,1577.8,345.39,580.07,681.38,0.0000,-3579.8,-6623.8,-299.55,-2717.9,-2550.5,-13692.,-1691.6,-1318.0,-5208.6,-2824.1,-5712.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1178.000000000,5759.5,1398.9,1546.5,1450.8,1801.3,1197.9,2651.6,494.73,1584.6,343.99,581.64,685.25,0.0000,-3573.9,-6615.3,-298.62,-2717.4,-2547.7,-13692.,-1690.2,-1314.7,-5207.1,-2823.6,-5711.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1179.000000000,5764.7,1397.3,1571.8,1451.6,1804.1,1216.4,2651.8,489.24,1598.6,346.78,574.55,682.71,0.0000,-3612.2,-6632.3,-301.91,-2717.2,-2573.4,-13693.,-1690.4,-1332.4,-5218.2,-2825.5,-5718.9,8594.9,3841.7,2942.9,2762.0,5354.2,1845.0,6613.5,1911.1,2921.7,872.08,1253.3,1509.7,0.0000,-8.7422,-9.0769,-1.3914,-8.3192,-5.4897,-33.686,-27.262,-2.7829,-24.464,-2.9693,-33.372
1180.000000000,5764.7,1393.1,1580.5,1456.9,1790.8,1200.3,2626.6,491.91,1606.1,345.01,573.00,683.84,0.0000,-3586.2,-6628.9,-301.16,-2717.0,-2554.6,-13693.,-1689.4,-1323.2,-5209.6,-2823.7,-5713.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1181.000000000,5725.0,1401.1,1583.7,1453.3,1791.0,1197.2,2606.0,490.56,1609.1,341.46,576.55,684.01,0.0000,-3578.6,-6622.2,-299.98,-2717.1,-2550.3,-13693.,-1688.6,-1318.7,-5206.7,-2822.9,-5711.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1182.000000000,5707.8,1401.2,1571.9,1451.7,1793.2,1190.2,2598.5,489.96,1591.8,341.66,580.73,684.70,0.0000,-3573.5,-6615.0,-298.95,-2717.2,-2547.3,-13693.,-1688.0,-1315.7,-5205.8,-2822.1,-5709.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1183.000000000,5686.9,1384.0,1573.1,1441.9,1794.4,1182.9,2592.0,487.46,1576.6,345.88,569.52,683.19,0.0000,-3568.7,-6608.5,-298.12,-2717.9,-2544.8,-13693.,-1687.6,-1313.2,-5206.0,-2820.8,-5709.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1184.000000000,5670.5,1392.2,1558.9,1439.7,1811.1,1204.0,2585.9,485.41,1579.2,344.11,568.79,680.87,0.0000,-3564.7,-6602.0,-297.45,-2718.8,-2542.4,-13692.,-1687.2,-1311.0,-5205.5,-2819.4,-5708.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1185.000000000,5585.8,1414.2,1565.4,1440.2,1805.6,1214.4,2561.1,477.91,1559.9,342.09,563.81,672.38,0.0000,-3561.5,-6597.0,-296.90,-2719.6,-2540.2,-13692.,-1687.0,-1308.7,-5204.8,-2817.8,-5707.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1186.000000000,5511.6,1435.2,1575.0,1445.9,1812.2,1208.2,2535.3,476.99,1545.9,342.45,558.98,659.41,0.0000,-3558.1,-6593.0,-296.43,-2720.2,-2538.1,-13691.,-1686.8,-1306.6,-5203.9,-2816.4,-5706.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1187.000000000,5495.6,1449.8,1582.4,1447.3,1819.3,1225.8,2545.7,478.52,1558.8,339.12,556.86,661.30,0.0000,-3598.8,-6612.0,-300.04,-2721.1,-2564.3,-13691.,-1686.8,-1324.4,-5214.2,-2817.8,-5713.6,1392.2,622.27,476.67,447.38,867.25,298.85,1071.2,309.56,473.24,141.26,203.01,244.53,0.0000,-1.4129,-1.4687,-0.22538,-1.3458,-0.88646,-5.4548,-4.4134,-0.45076,-3.9616,-0.48063,-5.4017
1188.000000000,5482.7,1423.5,1569.1,1434.5,1887.7,1208.3,2522.8,474.81,1549.4,341.69,562.62,663.71,0.0000,-3574.0,-6609.6,-299.51,-2721.9,-2546.2,-13690.,-1686.7,-1315.9,-5205.8,-2816.0,-5707.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1189.000000000,5488.4,1409.6,1556.5,1427.5,1877.3,1209.1,2507.2,476.37,1548.4,342.06,563.88,660.25,0.0000,-3566.7,-6603.1,-298.50,-2722.4,-2542.4,-13689.,-1686.5,-1311.7,-5203.4,-2815.7,-5705.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1190.000000000,5511.4,1425.2,1552.3,1424.8,1884.3,1202.3,2515.6,482.56,1540.9,340.04,567.32,657.75,0.0000,-3561.7,-6596.7,-297.64,-2722.3,-2539.7,-13688.,-1686.4,-1309.0,-5202.4,-2815.4,-5704.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1191.000000000,5513.5,1435.0,1551.6,1437.5,1878.4,1202.9,2540.6,478.46,1539.2,342.57,573.31,659.50,0.0000,-3557.2,-6591.1,-296.94,-2722.2,-2537.3,-13687.,-1686.3,-1306.8,-5201.6,-2814.9,-5704.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1192.000000000,5517.3,1442.3,1556.2,1431.9,1900.4,1197.5,2546.8,470.87,1545.0,342.09,566.49,666.47,0.0000,-3553.1,-6585.7,-296.37,-2722.1,-2535.3,-13687.,-1686.1,-1304.9,-5200.9,-2814.4,-5703.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1193.000000000,5479.9,1446.1,1547.1,1425.5,1880.2,1199.1,2555.0,472.67,1514.6,340.02,570.11,669.52,0.0000,-3549.3,-6580.7,-295.90,-2722.0,-2533.4,-13686.,-1686.0,-1303.3,-5200.4,-2813.7,-5702.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1194.000000000,5389.9,1437.3,1542.2,1432.4,1884.3,1198.9,2566.0,478.93,1498.7,337.93,569.07,662.61,0.0000,-3545.7,-6576.5,-295.49,-2722.0,-2531.5,-13685.,-1686.0,-1301.7,-5199.9,-2812.9,-5702.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1195.000000000,5353.8,1430.9,1550.8,1441.9,1882.1,1201.1,2579.4,483.01,1521.5,340.00,567.08,664.34,0.0000,-3542.4,-6572.5,-295.13,-2721.8,-2529.6,-13684.,-1685.9,-1300.3,-5199.6,-2812.0,-5701.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1196.000000000,5456.4,1425.1,1571.4,1424.6,1873.9,1200.5,2581.2,483.87,1523.4,339.61,572.00,660.76,0.0000,-3539.2,-6569.7,-294.80,-2721.6,-2527.8,-13683.,-1685.8,-1299.0,-5199.3,-2811.2,-5700.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1197.000000000,5448.8,1431.3,1593.1,1430.2,1863.2,1226.1,2567.0,484.75,1530.6,341.85,573.96,661.28,0.0000,-3579.5,-6590.5,-298.48,-2721.5,-2553.7,-13682.,-1686.1,-1316.6,-5210.5,-2812.6,-5708.4,2226.7,995.30,762.43,715.57,1387.2,478.01,1713.4,495.13,756.93,225.94,324.71,391.13,0.0000,-2.2528,-2.3451,-0.36049,-2.1498,-1.4120,-8.7227,-7.0534,-0.72097,-6.3341,-0.76842,-8.6304
1198.000000000,5438.1,1428.0,1581.6,1412.2,1884.0,1217.4,2573.1,484.21,1530.8,340.71,574.87,663.67,0.0000,-3555.1,-6590.0,-297.98,-2721.4,-2535.1,-13680.,-1685.9,-1309.1,-5202.5,-2810.2,-5702.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1199.000000000,5436.0,1440.4,1589.3,1413.2,1881.9,1227.4,2556.1,482.14,1536.0,343.20,576.27,667.01,0.0000,-3592.0,-6608.6,-300.97,-2721.4,-2558.9,-13679.,-1693.6,-1325.1,-5213.4,-2811.6,-5710.6,58026.,25937.,19868.,18647.,36148.,12456.,44649.,12903.,19725.,5887.7,8461.6,10192.,0.0000,-58.778,-61.143,-9.3939,-56.055,-36.807,-227.29,-183.78,-18.788,-165.05,-20.024,-224.85
1200.000000000,5436.6,1439.4,1586.7,1395.1,1910.2,1215.9,2536.9,478.95,1516.1,341.53,579.36,673.50,0.0000,-3566.1,-6605.6,-299.89,-2721.4,-2539.5,-13677.,-1691.6,-1315.5,-5205.4,-2809.3,-5705.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1201.000000000,5384.0,1432.8,1593.5,1371.0,1914.8,1215.8,2539.9,474.66,1500.8,342.30,578.94,681.90,0.0000,-3558.3,-6599.0,-298.45,-2721.3,-2535.1,-13676.,-1689.8,-1310.7,-5203.0,-2808.2,-5703.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1202.000000000,5372.8,1432.4,1598.2,1368.8,1919.3,1208.4,2523.6,470.60,1501.9,344.76,576.40,689.51,0.0000,-3552.6,-6592.5,-297.26,-2721.2,-2532.3,-13674.,-1688.5,-1307.4,-5201.5,-2807.3,-5702.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1203.000000000,5245.6,1443.9,1603.0,1384.3,1915.2,1212.9,2536.6,470.56,1506.8,343.12,576.99,692.50,0.0000,-3591.6,-6609.7,-300.34,-2721.1,-2557.9,-13674.,-1739.2,-1324.5,-5222.4,-2809.1,-5722.5,0.38506E+06,0.17211E+06,0.13184E+06,0.12374E+06,0.23988E+06,82660.,0.29629E+06,85621.,0.13089E+06,39070.,56151.,67637.,0.0000,-390.13,-405.84,-62.338,-372.02,-243.99,-1508.1,-1219.8,-124.68,-1095.1,-132.86,-1491.6
1204.000000000,5305.3,1568.9,1686.3,1380.0,1959.6,1335.3,2710.0,493.48,1510.3,362.57,615.57,739.51,0.0000,-3615.6,-6632.1,-303.55,-2723.0,-2574.1,-13679.,-1736.8,-1336.0,-5233.7,-2812.6,-5734.1,84674.,37848.,28992.,27210.,52748.,18177.,65154.,18828.,28783.,8591.5,12348.,14873.,0.0000,-86.274,-89.437,-13.708,-82.079,-54.204,-332.44,-268.53,-27.416,-240.97,-29.250,-328.51
1205.000000000,5311.5,1552.2,1734.1,1378.1,1958.9,1290.4,2635.0,486.32,1514.2,368.98,629.55,739.14,0.0000,-3635.2,-6655.1,-306.23,-2724.4,-2583.1,-13683.,-1723.3,-1345.1,-5239.6,-2816.1,-5736.3,2171.9,970.80,743.66,697.95,1353.0,466.24,1671.2,482.94,738.30,220.37,316.71,381.50,0.0000,-2.2204,-2.2964,-0.35161,-2.1092,-1.3962,-8.5330,-6.8912,-0.70322,-6.1829,-0.75056,-8.4322
1206.000000000,5364.2,1585.5,1713.8,1372.1,1969.7,1273.4,2617.3,484.47,1527.6,367.65,640.83,750.56,0.0000,-3652.4,-6672.3,-308.41,-2726.5,-2589.9,-13685.,-1712.9,-1352.9,-5239.7,-2819.6,-5734.9,2076.8,928.28,711.09,667.38,1293.7,445.82,1598.0,461.79,705.96,210.72,302.84,364.79,0.0000,-2.1287,-2.1979,-0.33621,-2.0195,-1.3383,-8.1615,-6.5916,-0.67242,-5.9134,-0.71782,-8.0668
1207.000000000,5353.0,1580.5,1704.4,1354.1,1940.7,1230.2,2612.6,494.62,1529.6,362.42,653.68,753.91,0.0000,-3622.0,-6664.8,-306.22,-2727.2,-2567.0,-13686.,-1705.0,-1337.6,-5226.7,-2820.9,-5724.1,509.77,227.86,174.54,163.82,317.56,109.43,392.25,113.35,173.29,51.724,74.336,89.542,0.0000,-0.52216,-0.53957,-0.82527E-01,-0.49541,-0.32782,-2.0030,-1.6182,-0.16505,-1.4516,-0.17619,-1.9804
1208.000000000,5248.7,1591.2,1719.3,1348.8,1944.9,1205.3,2599.8,501.79,1547.7,363.78,676.16,746.90,0.0000,-3611.2,-6654.4,-304.01,-2726.8,-2560.9,-13686.,-1699.5,-1330.5,-5221.1,-2823.8,-5718.4,1332.5,595.58,456.23,428.19,830.06,286.03,1025.3,296.28,452.94,135.20,194.30,234.05,0.0000,-1.3633,-1.4102,-0.21571,-1.2941,-0.85508,-5.2341,-4.2299,-0.43143,-3.7944,-0.46057,-5.1768
1209.000000000,5217.8,1597.4,1706.8,1338.8,1973.5,1185.7,2582.8,505.19,1539.6,362.23,678.29,749.16,0.0000,-3604.0,-6644.8,-302.31,-2725.5,-2556.7,-13686.,-1695.6,-1325.7,-5217.1,-2826.3,-5715.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1210.000000000,5213.8,1597.5,1713.6,1344.3,2028.9,1197.7,2600.3,513.62,1532.4,353.83,657.01,736.83,0.0000,-3643.4,-6657.8,-305.06,-2724.4,-2580.8,-13687.,-1693.7,-1343.3,-5225.5,-2828.5,-5720.4,6043.9,2701.5,2069.4,1942.2,3765.1,1297.4,4650.6,1343.9,2054.5,613.25,881.34,1061.6,0.0000,-6.1853,-6.3977,-0.97846,-5.8680,-3.8748,-23.733,-19.186,-1.9569,-17.211,-2.0891,-23.480
1211.000000000,5215.9,1561.3,1704.1,1334.0,2023.1,1189.5,2632.0,518.04,1539.3,353.98,645.87,725.53,0.0000,-3616.9,-6649.8,-303.92,-2723.2,-2560.3,-13687.,-1691.5,-1332.0,-5215.1,-2825.2,-5713.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1212.000000000,5207.1,1578.5,1695.1,1330.8,2035.5,1201.0,2657.2,522.51,1538.9,360.30,633.47,716.27,0.0000,-3608.2,-6638.9,-302.46,-2722.4,-2554.8,-13688.,-1690.0,-1326.1,-5211.8,-2822.8,-5710.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1213.000000000,5209.7,1584.6,1730.6,1325.3,2037.4,1214.8,2631.3,513.92,1541.0,363.79,623.26,723.59,0.0000,-3647.1,-6653.3,-305.26,-2721.9,-2579.1,-13689.,-1694.1,-1343.1,-5222.2,-2823.4,-5718.0,38107.,17033.,13048.,12246.,23739.,8180.4,29322.,8473.4,12954.,3866.6,5556.9,6693.6,0.0000,-38.991,-40.351,-6.1692,-36.981,-24.363,-149.56,-120.95,-12.338,-108.51,-13.165,-148.00
1214.000000000,5122.7,1565.7,1742.8,1298.8,2140.9,1191.2,2617.6,512.27,1526.2,366.10,618.76,724.54,0.0000,-3620.5,-6647.1,-304.12,-2721.6,-2559.0,-13689.,-1692.0,-1331.6,-5213.3,-2819.9,-5712.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1215.000000000,5142.8,1553.3,1723.6,1290.1,2179.3,1189.9,2620.3,514.57,1522.1,364.55,628.14,721.49,0.0000,-3611.2,-6638.1,-302.68,-2721.3,-2553.8,-13690.,-1690.4,-1325.6,-5210.0,-2818.1,-5710.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1216.000000000,5076.8,1533.6,1707.5,1301.8,2062.8,1198.5,2600.5,508.96,1517.6,364.17,631.19,726.80,0.0000,-3604.4,-6630.1,-301.49,-2721.1,-2550.3,-13690.,-1689.3,-1321.5,-5208.2,-2817.8,-5708.8,1128.1,504.24,386.26,362.52,702.76,242.17,868.04,250.84,383.48,114.46,164.50,198.15,0.0000,-1.1516,-1.1943,-0.18263,-1.0937,-0.71883,-4.4262,-3.5798,-0.36526,-3.2120,-0.38954,-4.3801
1217.000000000,5085.9,1514.7,1713.9,1317.6,1994.8,1189.5,2584.1,511.03,1514.2,365.14,629.45,731.14,0.0000,-3598.4,-6623.8,-300.54,-2720.7,-2547.2,-13690.,-1688.4,-1318.3,-5207.2,-2817.3,-5708.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1218.000000000,5082.9,1486.4,1739.3,1327.1,1968.5,1192.8,2569.5,509.03,1536.5,364.60,624.33,737.36,0.0000,-3637.1,-6640.8,-303.79,-2720.6,-2572.4,-13691.,-1687.9,-1336.7,-5217.7,-2819.4,-5715.5,1452.6,649.30,497.38,466.81,904.93,311.83,1117.8,323.00,493.80,147.39,211.83,255.16,0.0000,-1.4839,-1.5382,-0.23517,-1.4084,-0.92658,-5.6990,-4.6088,-0.47034,-4.1358,-0.50150,-5.6387
1219.000000000,5077.4,1478.9,1735.1,1332.4,1967.2,1169.5,2568.3,505.73,1528.1,360.80,621.30,739.27,0.0000,-3610.9,-6636.6,-302.96,-2720.5,-2553.0,-13691.,-1687.4,-1327.2,-5209.0,-2817.5,-5709.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1220.000000000,5059.5,1477.8,1736.9,1326.9,1953.4,1158.8,2584.9,504.82,1528.5,364.02,617.25,739.77,0.0000,-3602.4,-6628.2,-301.70,-2720.5,-2548.4,-13690.,-1687.0,-1322.4,-5207.0,-2816.4,-5707.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1221.000000000,5045.8,1473.6,1729.5,1314.1,1977.9,1157.6,2548.6,502.96,1533.3,365.29,608.37,739.43,0.0000,-3596.2,-6619.6,-300.61,-2720.9,-2545.5,-13690.,-1686.7,-1318.9,-5206.3,-2814.9,-5706.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1222.000000000,5020.1,1496.8,1737.7,1318.4,1965.0,1184.5,2546.3,501.27,1549.0,364.90,614.06,735.13,0.0000,-3591.2,-6611.8,-299.74,-2721.0,-2543.2,-13690.,-1686.4,-1316.0,-5205.4,-2813.9,-5705.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1223.000000000,5023.8,1506.6,1747.2,1325.5,1949.9,1182.5,2544.5,494.47,1539.1,364.62,607.91,726.58,0.0000,-3586.8,-6606.8,-299.04,-2720.8,-2540.8,-13689.,-1686.2,-1313.2,-5204.6,-2813.1,-5704.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1224.000000000,5226.4,1522.8,1752.5,1333.4,1928.6,1191.0,2531.3,495.66,1539.6,360.12,605.06,723.73,0.0000,-3582.6,-6602.4,-298.46,-2720.6,-2538.3,-13688.,-1686.1,-1310.8,-5203.5,-2812.2,-5703.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1225.000000000,5310.6,1525.9,1757.9,1345.7,1922.8,1220.8,2532.1,495.93,1550.8,358.19,604.19,732.59,0.0000,-3622.6,-6621.5,-301.96,-2720.5,-2564.4,-13689.,-1687.7,-1328.5,-5214.5,-2814.1,-5711.8,12455.,5567.1,4264.6,4002.4,7758.9,2673.7,9583.7,2769.4,4233.8,1263.7,1816.2,2187.7,0.0000,-12.694,-13.177,-2.0163,-12.061,-7.9283,-48.867,-39.494,-4.0327,-35.451,-4.2978,-48.311
1226.000000000,5353.0,1489.3,1731.9,1321.1,1910.7,1196.3,2511.8,493.93,1562.3,359.49,605.72,739.25,0.0000,-3596.7,-6618.6,-301.32,-2720.2,-2545.7,-13689.,-1687.2,-1319.5,-5206.1,-2812.3,-5706.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1227.000000000,5374.0,1475.4,1740.4,1317.9,1904.7,1180.5,2485.5,492.40,1561.1,356.84,611.70,741.79,0.0000,-3588.5,-6612.1,-300.19,-2719.6,-2541.3,-13689.,-1686.7,-1315.1,-5203.6,-2811.6,-5704.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1228.000000000,5314.7,1477.2,1746.2,1323.4,1896.9,1188.7,2458.2,490.14,1552.7,353.63,610.50,736.59,0.0000,-3582.5,-6605.5,-299.19,-2718.8,-2538.2,-13689.,-1686.4,-1312.1,-5202.2,-2810.8,-5703.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1229.000000000,5282.9,1496.9,1744.9,1333.8,1877.8,1222.1,2472.9,486.78,1552.9,351.52,610.20,737.46,0.0000,-3621.4,-6622.9,-302.39,-2718.1,-2563.6,-13690.,-1686.4,-1329.6,-5212.5,-2812.8,-5711.3,1597.5,714.07,547.00,513.38,995.20,342.94,1229.3,355.23,543.06,162.10,232.96,280.61,0.0000,-1.6277,-1.6899,-0.25863,-1.5466,-1.0159,-6.2679,-5.0639,-0.51726,-4.5463,-0.55115,-6.1937
1230.000000000,5247.1,1467.5,1737.5,1335.6,1873.9,1206.4,2462.6,485.84,1553.6,351.63,612.10,738.35,0.0000,-3595.5,-6620.3,-301.53,-2717.6,-2544.5,-13690.,-1686.1,-1320.5,-5203.7,-2810.8,-5705.7,146.02,65.270,49.999,46.925,90.967,31.347,112.36,32.470,49.638,14.816,21.294,25.649,0.0000,-0.14871,-0.15446,-0.23640E-01,-0.14134,-0.92735E-01,-0.57292,-0.46282,-0.47280E-01,-0.41554,-0.50375E-01,-0.56607
1231.000000000,5173.3,1460.4,1726.6,1335.1,1869.9,1232.5,2468.2,488.31,1575.6,351.86,616.59,737.90,0.0000,-3631.7,-6637.6,-304.27,-2717.2,-2567.9,-13691.,-1688.6,-1336.5,-5213.0,-2812.1,-5712.3,19940.,8912.7,6827.4,6407.7,12422.,4280.4,15343.,4433.8,6778.2,2023.2,2907.7,3502.5,0.0000,-20.343,-21.102,-3.2281,-19.312,-12.683,-78.234,-63.195,-6.4562,-56.740,-6.8792,-77.290
1232.000000000,5219.4,1457.1,1733.4,1342.0,1844.5,1229.9,2467.3,489.75,1580.7,350.98,613.72,739.51,0.0000,-3648.9,-6657.1,-307.01,-2717.0,-2576.1,-13691.,-1689.5,-1347.4,-5215.9,-2812.1,-5714.9,12461.,5569.8,4266.6,4004.4,7762.7,2675.0,9588.3,2770.8,4235.9,1264.4,1817.1,2188.8,0.0000,-12.739,-13.196,-2.0173,-12.080,-7.9350,-48.890,-39.490,-4.0346,-35.458,-4.2991,-48.296
1233.000000000,5118.3,1442.0,1689.7,1338.9,1777.8,1223.6,2469.3,490.05,1560.0,346.18,616.51,741.33,0.0000,-3618.4,-6651.5,-305.21,-2717.0,-2554.4,-13690.,-1688.5,-1334.0,-5205.3,-2809.2,-5707.7,367.67,164.34,125.89,118.15,229.04,78.926,282.91,81.753,124.98,37.305,53.614,64.581,0.0000,-0.37570,-0.38941,-0.59522E-01,-0.35634,-0.23373,-1.4425,-1.1651,-0.11904,-1.0461,-0.12684,-1.4248
1234.000000000,5244.3,1433.5,1668.0,1346.1,1826.2,1231.1,2469.7,485.10,1556.8,343.18,613.84,742.21,0.0000,-3652.5,-6664.8,-307.20,-2717.1,-2576.9,-13690.,-1693.9,-1348.8,-5214.7,-2810.3,-5714.9,46614.,20836.,15961.,14980.,29038.,10006.,35868.,10365.,15845.,4729.7,6797.4,8187.8,0.0000,-47.714,-49.397,-7.5464,-45.208,-29.674,-182.88,-147.71,-15.093,-132.63,-16.081,-180.63
1235.000000000,5244.2,1432.4,1680.3,1364.1,1871.4,1219.5,2459.8,484.59,1544.7,344.76,608.69,741.23,0.0000,-3668.0,-6680.2,-309.40,-2717.2,-2584.5,-13690.,-1708.0,-1358.4,-5220.6,-2810.6,-5721.6,0.12193E+06,54500.,41749.,39183.,75957.,26174.,93821.,27112.,41448.,12372.,17780.,21417.,0.0000,-125.05,-129.30,-19.739,-118.37,-77.700,-478.35,-386.40,-39.479,-346.92,-42.066,-472.45
1236.000000000,5217.8,1427.5,1695.0,1381.8,1873.8,1221.7,2467.1,486.50,1543.2,337.91,609.22,730.86,0.0000,-3680.7,-6694.9,-311.28,-2717.4,-2590.2,-13690.,-1705.4,-1365.9,-5223.1,-2810.5,-5724.9,24398.,10906.,8354.0,7840.5,15199.,5237.5,18774.,5425.2,8293.8,2475.6,3557.9,4285.6,0.0000,-25.072,-25.895,-3.9499,-23.706,-15.561,-95.725,-77.323,-7.8998,-69.418,-8.4176,-94.535
1237.000000000,5214.8,1434.6,1737.8,1388.6,1886.5,1199.2,2497.3,494.33,1525.2,336.70,609.07,737.50,0.0000,-3647.8,-6684.3,-308.81,-2717.6,-2568.7,-13690.,-1699.9,-1349.0,-5211.3,-2808.0,-5717.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1238.000000000,5230.2,1444.8,1744.1,1395.8,1882.8,1179.8,2501.4,494.65,1511.0,338.86,622.74,732.43,0.0000,-3637.4,-6671.7,-306.32,-2717.5,-2563.7,-13691.,-1695.7,-1340.5,-5206.8,-2807.2,-5713.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1239.000000000,5216.3,1423.5,1741.0,1405.2,1873.6,1157.4,2465.9,493.28,1517.8,339.04,621.38,735.58,0.0000,-3628.9,-6659.4,-304.38,-2717.1,-2559.7,-13692.,-1692.6,-1334.6,-5204.8,-2806.5,-5710.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1240.000000000,5251.9,1433.9,1740.2,1412.4,1880.0,1164.0,2477.2,495.83,1519.4,338.45,622.67,734.85,0.0000,-3621.2,-6647.2,-302.92,-2716.7,-2556.2,-13692.,-1690.4,-1330.0,-5203.0,-2806.0,-5708.6,5.2831,2.3614,1.8089,1.6977,3.2911,1.1341,4.0652,1.1747,1.7959,0.53605,0.77040,0.92798,0.0000,-0.54170E-02,-0.56075E-02,-0.85528E-03,-0.51279E-02,-0.33664E-02,-0.20747E-01,-0.16749E-01,-0.17106E-02,-0.15035E-01,-0.18229E-02,-0.20482E-01
1241.000000000,5245.4,1431.5,1747.8,1417.4,1877.5,1166.9,2500.6,495.29,1515.0,337.74,622.08,736.35,0.0000,-3614.4,-6636.8,-301.80,-2716.5,-2552.8,-13692.,-1688.9,-1326.1,-5201.5,-2805.9,-5707.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1242.000000000,5242.0,1435.0,1737.3,1427.3,1881.9,1161.9,2499.0,492.99,1517.6,339.51,618.09,731.55,0.0000,-3607.9,-6627.7,-300.92,-2715.8,-2549.3,-13692.,-1687.8,-1322.7,-5200.2,-2805.5,-5706.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1243.000000000,5208.2,1448.1,1716.8,1441.6,1886.6,1161.9,2499.5,493.64,1522.8,338.97,619.69,735.61,0.0000,-3601.8,-6619.4,-300.21,-2715.1,-2546.0,-13693.,-1687.2,-1319.7,-5199.3,-2805.0,-5705.3,1061.0,474.24,363.28,340.95,660.95,227.76,816.39,235.92,360.66,107.65,154.72,186.36,0.0000,-1.0844,-1.1248,-0.17176,-1.0284,-0.67425,-4.1663,-3.3633,-0.34353,-3.0193,-0.36601,-4.1129
1244.000000000,5205.9,1434.2,1701.6,1433.7,1900.4,1163.6,2519.4,492.55,1529.2,337.28,627.73,732.76,0.0000,-3596.1,-6612.5,-299.61,-2714.3,-2542.8,-13693.,-1686.6,-1317.1,-5198.5,-2804.6,-5704.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1245.000000000,5200.7,1429.1,1707.9,1431.6,1899.2,1160.6,2505.2,496.72,1523.0,338.60,632.19,734.92,0.0000,-3590.5,-6607.6,-299.08,-2713.5,-2539.6,-13694.,-1686.1,-1314.8,-5197.9,-2804.4,-5703.9,8.8141,3.9397,3.0179,2.8324,5.4908,1.8921,6.7822,1.9599,2.9962,0.89432,1.2853,1.5482,0.0000,-0.89907E-02,-0.93357E-02,-0.14269E-02,-0.85369E-02,-0.55899E-02,-0.34608E-01,-0.27936E-01,-0.28538E-02,-0.25082E-01,-0.30405E-02,-0.34161E-01
1246.000000000,5176.2,1439.6,1716.7,1428.8,1909.3,1181.4,2496.6,498.36,1527.3,338.75,628.90,735.51,0.0000,-3629.1,-6626.0,-302.62,-2712.6,-2564.7,-13695.,-1686.6,-1333.0,-5208.7,-2806.8,-5711.5,5476.8,2448.0,1875.2,1760.0,3411.8,1175.7,4214.2,1217.8,1861.7,555.70,798.64,962.01,0.0000,-5.5951,-5.8021,-0.88664,-5.3072,-3.4789,-21.504,-17.358,-1.7733,-15.585,-1.8893,-21.224
1247.000000000,5128.8,1443.3,1724.1,1402.3,1878.0,1183.7,2508.3,499.28,1520.9,337.45,634.02,731.69,0.0000,-3602.5,-6623.5,-301.99,-2711.6,-2545.3,-13694.,-1686.2,-1323.8,-5200.2,-2805.6,-5705.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1248.000000000,5099.3,1446.0,1722.5,1402.7,1903.2,1190.2,2503.3,504.57,1527.1,339.06,633.50,729.10,0.0000,-3638.2,-6641.0,-304.88,-2710.7,-2568.3,-13694.,-1687.8,-1340.0,-5209.2,-2807.8,-5712.6,13916.,6220.3,4764.9,4472.1,8669.3,2987.4,10708.,3094.4,4730.6,1412.0,2029.3,2444.4,0.0000,-14.232,-14.747,-2.2529,-13.491,-8.8389,-54.638,-44.099,-4.5059,-39.598,-4.8006,-53.920
1249.000000000,5099.8,1447.8,1700.9,1382.8,1918.8,1193.5,2515.5,505.21,1529.1,339.57,626.12,726.35,0.0000,-3655.3,-6659.6,-307.71,-2710.1,-2576.1,-13694.,-1720.5,-1350.8,-5218.5,-2808.5,-5723.7,0.25008E+06,0.11178E+06,85626.,80363.,0.15579E+06,53683.,0.19243E+06,55606.,85009.,25374.,36467.,43926.,0.0000,-256.26,-265.16,-40.485,-242.66,-158.99,-981.85,-792.66,-80.970,-711.57,-86.269,-968.89
1250.000000000,5233.7,1469.9,1705.1,1364.9,1884.3,1204.7,2526.3,511.35,1527.0,343.85,621.97,738.83,0.0000,-3669.4,-6676.9,-310.02,-2709.8,-2582.9,-13695.,-1718.9,-1359.4,-5224.0,-2808.7,-5730.8,54884.,24532.,18792.,17637.,34190.,11782.,42231.,12204.,18657.,5568.8,8003.4,9640.5,0.0000,-56.370,-58.253,-8.8852,-53.326,-34.955,-215.59,-174.01,-17.770,-156.18,-18.933,-212.71
1251.000000000,5209.7,1558.2,1754.3,1362.0,1879.4,1267.7,2599.2,520.31,1519.1,351.38,642.74,753.73,0.0000,-3686.3,-6695.0,-311.93,-2710.4,-2591.8,-13698.,-1710.5,-1366.7,-5225.7,-2810.5,-5732.6,5055.9,2259.9,1731.1,1624.7,3149.6,1085.3,3890.4,1124.2,1718.7,513.00,737.27,888.08,0.0000,-5.2144,-5.3733,-0.81851,-4.9229,-3.2358,-19.880,-16.037,-1.6370,-14.392,-1.7455,-19.606
1252.000000000,5253.1,1535.1,1730.1,1362.6,1875.7,1234.1,2556.2,507.22,1497.2,351.89,634.31,758.00,0.0000,-3655.1,-6686.1,-309.47,-2710.4,-2569.7,-13700.,-1703.3,-1349.9,-5214.7,-2808.9,-5723.4,2.1282,0.95125,0.72869,0.68390,1.3258,0.45685,1.6376,0.47322,0.72343,0.21594,0.31034,0.37382,0.0000,-0.21943E-02,-0.22623E-02,-0.34453E-03,-0.20715E-02,-0.13612E-02,-0.83707E-02,-0.67518E-02,-0.68906E-03,-0.60586E-02,-0.73468E-03,-0.82553E-02
1253.000000000,5256.7,1545.4,1718.9,1371.2,1878.5,1213.9,2540.0,496.89,1492.8,350.84,634.63,756.25,0.0000,-3644.5,-6673.0,-306.95,-2710.6,-2563.5,-13701.,-1697.9,-1341.6,-5210.0,-2809.0,-5718.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1254.000000000,5252.4,1548.7,1705.9,1386.3,1870.5,1194.7,2537.4,493.95,1511.9,350.36,629.83,759.04,0.0000,-3636.4,-6660.0,-304.99,-2710.2,-2559.0,-13701.,-1694.1,-1335.9,-5206.8,-2809.3,-5715.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1255.000000000,5310.8,1533.1,1722.4,1387.2,1892.1,1199.3,2562.9,505.17,1516.3,349.10,643.20,756.21,0.0000,-3629.1,-6650.0,-303.55,-2709.5,-2555.2,-13702.,-1691.5,-1331.6,-5204.5,-2810.1,-5713.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1256.000000000,5313.0,1544.9,1727.6,1399.5,1880.4,1193.3,2559.1,508.64,1513.1,345.10,657.04,759.59,0.0000,-3622.6,-6641.1,-302.46,-2708.6,-2551.9,-13703.,-1689.7,-1328.0,-5202.3,-2811.5,-5711.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1257.000000000,5319.0,1518.4,1720.8,1396.3,1893.5,1199.4,2551.9,514.35,1510.7,344.05,655.53,759.38,0.0000,-3617.2,-6632.9,-301.61,-2707.6,-2548.6,-13704.,-1688.4,-1324.9,-5200.5,-2812.0,-5710.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1258.000000000,5344.0,1519.8,1705.1,1408.9,1887.0,1197.5,2576.6,522.43,1513.4,339.92,648.97,746.12,0.0000,-3612.2,-6624.7,-300.90,-2706.7,-2545.5,-13705.,-1687.5,-1322.1,-5198.7,-2811.4,-5709.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1259.000000000,5376.0,1516.0,1678.3,1413.6,1892.3,1192.7,2591.1,518.23,1518.7,343.72,644.49,726.03,0.0000,-3607.3,-6617.3,-300.29,-2705.9,-2542.3,-13706.,-1686.9,-1319.5,-5197.4,-2810.2,-5708.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1260.000000000,5378.5,1536.8,1679.2,1425.2,1908.1,1204.6,2588.4,509.52,1522.2,347.62,640.82,715.34,0.0000,-3646.8,-6634.3,-303.77,-2705.1,-2567.0,-13708.,-1686.8,-1337.8,-5208.0,-2811.4,-5716.0,2614.2,1168.5,895.11,840.09,1628.5,561.19,2011.6,581.29,888.65,265.25,381.21,459.19,0.0000,-2.6789,-2.7717,-0.42322,-2.5362,-1.6598,-10.273,-8.2921,-0.84644,-7.4419,-0.90188,-10.137
1261.000000000,5453.5,1508.3,1681.9,1433.7,1904.3,1190.4,2568.9,503.26,1507.0,348.31,631.50,718.34,0.0000,-3620.8,-6630.7,-303.08,-2704.5,-2547.1,-13708.,-1686.4,-1328.1,-5199.4,-2808.5,-5710.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1262.000000000,5478.2,1491.2,1680.0,1437.0,1929.4,1186.7,2554.9,502.00,1503.0,344.99,629.30,715.00,0.0000,-3612.2,-6623.6,-301.90,-2704.1,-2541.9,-13709.,-1686.0,-1323.3,-5196.7,-2807.0,-5708.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1263.000000000,5506.7,1475.4,1668.0,1440.9,1931.1,1199.1,2544.6,494.05,1503.2,344.35,634.63,713.91,0.0000,-3605.7,-6616.1,-300.85,-2703.8,-2538.5,-13708.,-1685.8,-1320.0,-5195.4,-2806.6,-5707.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1264.000000000,5521.7,1459.2,1686.1,1444.0,1919.7,1193.4,2546.8,485.55,1500.2,344.70,630.00,721.10,0.0000,-3599.9,-6611.0,-299.97,-2703.5,-2535.6,-13708.,-1685.6,-1317.2,-5195.1,-2806.3,-5707.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1265.000000000,5585.6,1431.3,1682.8,1440.2,1843.4,1192.9,2533.6,486.31,1502.4,340.98,627.08,716.29,0.0000,-3594.5,-6606.8,-299.23,-2703.2,-2532.8,-13706.,-1685.4,-1315.3,-5194.6,-2805.4,-5707.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1266.000000000,5677.3,1441.8,1687.1,1434.8,1819.9,1193.9,2554.4,483.77,1497.5,335.92,624.35,708.31,0.0000,-3589.8,-6602.3,-298.62,-2703.0,-2530.3,-13705.,-1685.2,-1313.4,-5194.0,-2804.5,-5706.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1267.000000000,5769.0,1433.0,1678.5,1431.0,1822.6,1218.3,2579.5,481.51,1509.3,337.91,629.63,715.03,0.0000,-3629.2,-6621.6,-302.10,-2702.9,-2555.9,-13705.,-1692.6,-1331.5,-5207.1,-2806.3,-5716.3,55308.,24722.,18938.,17774.,34455.,11873.,42558.,12298.,18801.,5611.9,8065.3,9715.0,0.0000,-56.484,-58.554,-8.9539,-53.580,-34.988,-217.24,-175.33,-17.908,-157.40,-19.066,-214.27
1268.000000000,5821.4,1431.7,1646.6,1434.5,1860.6,1216.1,2555.6,482.52,1509.0,340.93,628.38,713.45,0.0000,-3603.3,-6619.8,-301.44,-2703.3,-2537.0,-13704.,-1690.7,-1322.6,-5199.9,-2804.1,-5711.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1269.000000000,5798.4,1437.5,1639.8,1429.5,1862.9,1230.7,2539.3,483.60,1512.2,340.78,626.18,710.57,0.0000,-3595.5,-6614.4,-300.30,-2703.6,-2532.8,-13704.,-1689.0,-1318.2,-5197.6,-2802.8,-5710.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1270.000000000,5926.4,1426.0,1650.1,1423.5,1870.1,1212.4,2543.4,481.16,1485.7,337.45,627.96,699.73,0.0000,-3590.1,-6609.9,-299.28,-2703.7,-2530.1,-13703.,-1687.8,-1315.1,-5196.0,-2801.7,-5708.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1271.000000000,5922.3,1407.2,1646.8,1418.7,1871.5,1211.8,2550.2,479.45,1458.3,335.95,624.84,691.89,0.0000,-3585.1,-6605.3,-298.46,-2704.1,-2527.8,-13702.,-1686.9,-1312.6,-5194.9,-2800.7,-5707.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1272.000000000,5973.1,1391.3,1641.8,1423.4,1864.6,1209.8,2552.9,479.64,1456.5,335.97,625.91,685.57,0.0000,-3580.4,-6600.7,-297.77,-2704.6,-2526.0,-13701.,-1686.2,-1310.4,-5193.7,-2800.0,-5706.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1273.000000000,6135.5,1392.9,1628.9,1438.7,1858.9,1214.5,2541.0,480.51,1440.6,338.30,623.20,683.06,0.0000,-3620.0,-6619.4,-301.21,-2704.8,-2552.0,-13701.,-1692.9,-1328.1,-5205.6,-2802.1,-5715.8,53345.,23844.,18265.,17143.,33232.,11451.,41047.,11862.,18134.,5412.7,7778.9,9370.1,0.0000,-54.370,-56.413,-8.6361,-51.633,-33.683,-209.45,-169.04,-17.272,-151.78,-18.381,-206.50
1274.000000000,6221.5,1381.6,1625.5,1444.9,1853.3,1224.8,2579.4,485.32,1460.4,340.05,623.15,686.31,0.0000,-3638.5,-6639.6,-304.55,-2705.0,-2561.1,-13701.,-1747.0,-1340.1,-5220.9,-2802.7,-5733.8,0.41833E+06,0.18699E+06,0.14324E+06,0.13443E+06,0.26060E+06,89802.,0.32189E+06,93019.,0.14220E+06,42446.,61002.,73480.,0.0000,-427.27,-442.68,-67.724,-405.20,-264.51,-1642.6,-1326.3,-135.45,-1190.2,-144.15,-1619.5
1275.000000000,6200.4,1611.7,1760.5,1446.8,1911.1,1431.1,2902.2,514.34,1471.2,384.83,692.20,774.91,0.0000,-3663.8,-6666.4,-307.42,-2708.6,-2578.9,-13711.,-1733.1,-1349.8,-5232.1,-2808.5,-5742.5,14788.,6610.1,5063.5,4752.3,9212.5,3174.6,11379.,3288.3,5027.0,1500.5,2156.5,2597.6,0.0000,-15.232,-15.692,-2.3941,-14.397,-9.4887,-58.267,-46.952,-4.7882,-42.115,-5.1061,-57.376
1276.000000000,5955.8,1600.1,1742.8,1437.6,2068.0,1297.1,2702.4,492.76,1472.7,380.97,685.20,758.59,0.0000,-3683.2,-6686.2,-309.75,-2711.7,-2585.4,-13715.,-1720.6,-1358.0,-5237.3,-2813.4,-5744.0,4698.0,2099.9,1608.6,1509.7,2926.7,1008.5,3615.0,1044.6,1597.0,476.68,685.08,825.21,0.0000,-4.8505,-4.9881,-0.76057,-4.5797,-3.0215,-18.514,-14.922,-1.5211,-13.382,-1.6223,-18.237
1277.000000000,5936.1,1579.4,1698.6,1433.2,2055.0,1232.2,2652.5,499.68,1481.8,365.72,696.01,759.68,0.0000,-3652.8,-6678.5,-307.70,-2712.5,-2562.0,-13715.,-1710.4,-1343.0,-5224.2,-2815.3,-5734.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1278.000000000,5963.5,1584.3,1717.2,1417.9,2025.6,1195.0,2625.8,508.29,1487.5,364.25,726.38,738.18,0.0000,-3641.5,-6670.1,-305.59,-2711.7,-2555.4,-13716.,-1703.0,-1335.8,-5217.7,-2818.8,-5728.2,334.70,149.60,114.60,107.56,208.50,71.849,257.54,74.423,113.77,33.960,48.807,58.791,0.0000,-0.34468,-0.35519,-0.54185E-01,-0.32575,-0.21420,-1.3179,-1.0633,-0.10837,-0.95347,-0.11557,-1.2995
1279.000000000,6078.4,1558.7,1674.2,1425.1,2061.9,1180.6,2587.5,500.58,1475.0,362.99,703.73,733.30,0.0000,-3634.3,-6658.4,-303.94,-2710.7,-2550.5,-13715.,-1697.8,-1331.0,-5212.8,-2819.8,-5724.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1280.000000000,6144.9,1545.1,1682.9,1458.9,2069.7,1193.9,2644.6,522.04,1500.4,361.06,685.08,717.32,0.0000,-3628.3,-6648.5,-302.70,-2709.7,-2546.6,-13715.,-1694.1,-1327.2,-5208.5,-2818.6,-5721.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1281.000000000,6143.4,1556.2,1694.5,1472.9,2090.8,1229.0,2635.9,514.09,1510.8,367.13,678.88,715.40,0.0000,-3622.7,-6641.0,-301.76,-2708.4,-2543.3,-13715.,-1691.6,-1324.0,-5205.8,-2817.3,-5718.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1282.000000000,6258.3,1554.9,1719.9,1488.0,2103.7,1239.8,2622.7,508.31,1506.8,368.59,670.29,727.59,0.0000,-3618.2,-6635.1,-301.00,-2707.3,-2540.1,-13715.,-1689.9,-1321.2,-5203.7,-2815.5,-5717.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1283.000000000,6380.3,1538.4,1741.6,1488.3,2154.3,1212.3,2600.0,502.54,1512.4,374.65,643.77,738.22,0.0000,-3613.8,-6628.7,-300.36,-2706.5,-2537.0,-13715.,-1688.7,-1318.7,-5202.1,-2813.2,-5716.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1284.000000000,6298.5,1556.7,1732.1,1485.9,2186.9,1218.8,2608.1,496.83,1525.5,375.37,635.72,736.35,0.0000,-3609.1,-6621.0,-299.81,-2706.1,-2534.0,-13715.,-1687.8,-1316.4,-5200.8,-2811.0,-5715.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1285.000000000,6410.7,1545.0,1753.3,1490.5,2198.9,1224.3,2601.6,494.03,1525.9,382.41,641.98,746.33,0.0000,-3603.8,-6615.7,-299.32,-2705.8,-2531.4,-13715.,-1687.2,-1314.4,-5200.4,-2810.1,-5715.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1286.000000000,6395.3,1538.5,1793.6,1485.4,2199.6,1213.6,2574.5,495.35,1540.3,380.55,643.16,757.27,0.0000,-3598.6,-6612.0,-298.87,-2705.6,-2528.8,-13714.,-1686.8,-1313.2,-5200.2,-2809.5,-5715.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1287.000000000,6342.8,1512.0,1801.5,1478.4,2233.5,1202.3,2573.3,492.93,1539.4,375.80,643.46,757.48,0.0000,-3594.5,-6608.8,-298.45,-2705.6,-2526.3,-13714.,-1686.5,-1312.1,-5199.8,-2808.9,-5714.9,488.17,218.20,167.15,156.87,304.11,104.79,375.63,108.55,165.94,49.532,71.186,85.748,0.0000,-0.49784,-0.51647,-0.79030E-01,-0.47317,-0.30929,-1.9178,-1.5499,-0.15806,-1.3903,-0.16829,-1.8935
1288.000000000,6466.8,1507.3,1783.2,1477.5,2369.0,1197.6,2585.4,490.36,1545.1,381.42,641.00,747.97,0.0000,-3589.6,-6604.9,-298.06,-2706.5,-2524.1,-13714.,-1686.3,-1310.8,-5200.4,-2808.4,-5714.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1289.000000000,6591.2,1526.6,1782.5,1473.7,2320.9,1211.6,2584.1,487.57,1583.6,380.52,643.19,741.51,0.0000,-3585.6,-6601.9,-297.71,-2707.5,-2522.2,-13714.,-1686.0,-1309.6,-5200.4,-2808.0,-5714.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1290.000000000,6695.2,1528.1,1806.0,1474.9,2301.3,1210.4,2583.8,485.79,1582.5,381.34,628.69,735.76,0.0000,-3582.4,-6601.0,-297.37,-2708.4,-2520.3,-13714.,-1685.9,-1308.3,-5200.1,-2806.5,-5713.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1291.000000000,6872.2,1515.5,1793.2,1460.2,2328.8,1235.9,2581.9,482.05,1581.1,380.55,624.34,729.06,0.0000,-3579.5,-6598.4,-297.06,-2710.2,-2518.9,-13715.,-1685.7,-1306.9,-5199.0,-2805.0,-5712.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1292.000000000,7000.9,1503.3,1773.2,1450.3,2339.3,1255.2,2568.2,475.24,1611.9,386.21,626.72,722.13,0.0000,-3575.9,-6595.6,-296.75,-2711.7,-2517.6,-13715.,-1685.6,-1305.0,-5198.3,-2804.2,-5712.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1293.000000000,6799.6,1502.0,1771.7,1446.8,2330.2,1262.8,2539.0,476.12,1608.9,382.63,629.43,724.61,0.0000,-3572.2,-6592.7,-296.47,-2712.8,-2516.1,-13715.,-1685.5,-1303.5,-5196.9,-2803.6,-5711.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1294.000000000,6817.1,1529.7,1794.6,1432.9,2315.8,1256.5,2571.5,471.84,1583.9,376.88,630.07,731.02,0.0000,-3568.5,-6589.8,-296.20,-2713.1,-2514.4,-13715.,-1685.4,-1302.3,-5195.5,-2803.1,-5711.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1295.000000000,6844.2,1532.9,1655.7,1408.9,2322.5,1247.4,2568.6,472.42,1581.9,375.86,634.47,736.50,0.0000,-3564.2,-6585.2,-295.93,-2713.3,-2512.5,-13715.,-1685.4,-1301.4,-5194.7,-2802.4,-5711.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1296.000000000,6839.1,1532.8,1579.3,1414.5,2305.7,1235.7,2563.5,472.44,1609.6,375.98,636.64,730.70,0.0000,-3560.0,-6580.6,-295.68,-2713.0,-2510.5,-13716.,-1685.3,-1300.6,-5194.1,-2801.7,-5711.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1297.000000000,6730.9,1550.9,1593.3,1436.1,2317.6,1211.0,2552.7,474.17,1629.0,376.88,638.57,731.83,0.0000,-3556.0,-6578.0,-295.42,-2712.6,-2508.2,-13716.,-1685.2,-1299.9,-5193.5,-2800.6,-5711.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1298.000000000,6739.7,1548.1,1605.9,1446.9,2298.8,1232.5,2543.0,476.36,1633.1,375.09,642.96,735.97,0.0000,-3552.2,-6577.1,-295.16,-2712.4,-2506.2,-13715.,-1685.2,-1299.3,-5193.0,-2799.6,-5711.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1299.000000000,6671.0,1544.0,1627.9,1447.9,2294.5,1231.5,2471.4,480.15,1633.4,375.21,645.95,740.48,0.0000,-3548.5,-6576.0,-294.90,-2712.3,-2504.3,-13714.,-1685.1,-1298.5,-5193.0,-2798.6,-5710.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1300.000000000,6598.7,1521.9,1645.2,1453.5,2250.8,1214.3,2477.2,476.91,1633.1,379.57,642.87,745.05,0.0000,-3545.0,-6574.4,-294.64,-2712.2,-2502.6,-13713.,-1685.0,-1297.7,-5193.0,-2797.8,-5710.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1301.000000000,6526.5,1521.0,1658.6,1472.9,2317.0,1185.3,2475.1,471.87,1654.6,380.58,636.07,744.57,0.0000,-3541.6,-6572.7,-294.39,-2712.0,-2500.9,-13712.,-1685.0,-1296.8,-5192.8,-2797.0,-5710.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1302.000000000,6466.9,1524.2,1677.6,1485.1,2373.7,1183.9,2478.6,473.62,1682.1,379.90,631.02,750.69,0.0000,-3538.2,-6569.5,-294.14,-2711.8,-2499.2,-13710.,-1684.9,-1295.8,-5192.6,-2796.3,-5709.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1303.000000000,6450.7,1513.4,1675.0,1496.3,2337.6,1191.1,2458.3,466.11,1708.9,380.85,620.34,753.67,0.0000,-3578.4,-6588.8,-297.90,-2711.9,-2525.3,-13710.,-1685.1,-1312.5,-5203.8,-2798.2,-5717.8,1387.8,620.31,475.17,445.96,864.52,297.91,1067.8,308.58,471.74,140.81,202.37,243.76,0.0000,-1.4034,-1.4613,-0.22467,-1.3413,-0.87536,-5.4425,-4.3990,-0.44933,-3.9494,-0.47801,-5.3702
1304.000000000,6461.9,1500.3,1657.2,1496.5,2302.9,1200.8,2499.7,459.96,1738.3,381.45,620.75,746.86,0.0000,-3597.5,-6610.7,-301.49,-2711.9,-2534.7,-13710.,-1690.9,-1324.8,-5207.9,-2798.7,-5721.9,43539.,19461.,14908.,13991.,27123.,9346.4,33502.,9681.2,14800.,4417.7,6349.0,7647.7,0.0000,-44.104,-45.875,-7.0486,-42.111,-27.503,-170.73,-138.01,-14.097,-123.90,-14.997,-168.46
1305.000000000,6488.0,1517.0,1657.4,1501.3,2307.5,1216.9,2525.6,459.82,1726.2,382.54,620.53,745.60,0.0000,-3613.0,-6631.0,-304.38,-2712.0,-2541.9,-13711.,-1690.0,-1335.0,-5209.5,-2798.8,-5724.0,4022.2,1797.9,1377.2,1292.6,2505.7,863.44,3095.0,894.37,1367.3,408.12,586.53,706.51,0.0000,-4.0834,-4.2413,-0.65116,-3.8936,-2.5435,-15.771,-12.748,-1.3023,-11.446,-1.3855,-15.561
1306.000000000,6540.8,1493.5,1620.2,1509.0,2309.1,1201.6,2493.9,460.47,1718.9,382.47,621.66,737.69,0.0000,-3582.9,-6626.0,-302.62,-2712.0,-2520.3,-13711.,-1688.6,-1323.1,-5198.5,-2796.2,-5716.8,23.740,10.611,8.1286,7.6290,14.789,5.0962,18.267,5.2788,8.0700,2.4088,3.4619,4.1700,0.0000,-0.24094E-01,-0.25039E-01,-0.38433E-02,-0.22977E-01,-0.14987E-01,-0.93073E-01,-0.75237E-01,-0.76866E-02,-0.67554E-01,-0.81766E-02,-0.91832E-01
1307.000000000,6716.6,1470.1,1594.9,1536.6,2301.7,1242.2,2500.9,457.45,1711.1,378.28,627.34,731.78,0.0000,-3617.3,-6640.5,-304.60,-2712.0,-2542.8,-13712.,-1687.8,-1338.1,-5206.0,-2797.4,-5722.1,1816.7,812.04,622.05,583.81,1131.7,389.99,1397.9,403.96,617.56,184.33,264.92,319.11,0.0000,-1.8474,-1.9171,-0.29411,-1.7594,-1.1485,-7.1217,-5.7571,-0.58822,-5.1695,-0.62572,-7.0267
1308.000000000,6755.2,1488.0,1570.8,1534.8,2228.1,1251.4,2534.5,456.78,1714.4,373.60,633.62,728.20,0.0000,-3588.9,-6633.7,-302.77,-2711.9,-2522.8,-13711.,-1686.9,-1327.1,-5196.1,-2795.0,-5715.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1309.000000000,6766.6,1466.2,1569.5,1550.8,2201.8,1269.7,2523.1,464.23,1695.6,367.17,631.56,730.32,0.0000,-3579.2,-6624.2,-300.80,-2711.6,-2517.8,-13709.,-1686.2,-1321.5,-5192.8,-2793.8,-5712.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1310.000000000,6671.9,1426.6,1574.1,1540.7,2178.9,1279.3,2544.1,463.68,1701.5,367.13,628.75,726.38,0.0000,-3572.2,-6615.2,-299.22,-2711.3,-2514.6,-13707.,-1685.7,-1317.7,-5191.4,-2792.7,-5711.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1311.000000000,6605.7,1435.3,1546.1,1530.0,2193.3,1278.1,2544.6,457.25,1698.9,363.48,636.44,720.89,0.0000,-3566.0,-6607.7,-298.01,-2711.6,-2512.0,-13705.,-1685.3,-1314.4,-5190.6,-2791.7,-5709.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1312.000000000,6601.6,1474.7,1549.2,1563.4,2219.1,1231.0,2539.4,459.55,1713.7,363.22,644.22,710.78,0.0000,-3560.3,-6600.8,-297.06,-2711.8,-2509.6,-13703.,-1685.1,-1311.6,-5189.8,-2790.8,-5708.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1313.000000000,6582.3,1427.5,1561.2,1588.0,2221.1,1212.2,2582.2,460.55,1696.3,362.08,646.31,713.28,0.0000,-3555.1,-6594.6,-296.29,-2711.9,-2507.3,-13701.,-1684.8,-1309.2,-5189.2,-2790.0,-5708.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1314.000000000,6570.2,1435.2,1557.1,1580.8,2201.0,1206.4,2601.6,461.46,1685.3,358.38,642.91,709.14,0.0000,-3550.3,-6589.0,-295.65,-2711.9,-2505.2,-13700.,-1684.7,-1307.1,-5188.8,-2789.2,-5707.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1315.000000000,6494.4,1448.0,1550.4,1585.7,2208.4,1231.8,2562.4,460.63,1687.6,356.72,649.24,721.09,0.0000,-3545.8,-6585.4,-295.09,-2711.8,-2503.2,-13698.,-1684.5,-1305.2,-5188.6,-2788.5,-5706.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1316.000000000,6480.1,1462.3,1560.8,1595.7,2189.3,1241.3,2573.9,461.49,1674.9,358.91,643.07,728.42,0.0000,-3541.4,-6582.3,-294.59,-2710.9,-2501.3,-13696.,-1684.4,-1303.3,-5188.0,-2787.8,-5705.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1317.000000000,6523.9,1432.8,1559.3,1572.6,2126.7,1251.7,2550.0,469.18,1677.5,358.67,639.25,733.40,0.0000,-3537.5,-6579.2,-294.13,-2709.8,-2499.6,-13694.,-1684.3,-1301.6,-5187.4,-2787.1,-5704.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1318.000000000,6464.7,1430.1,1543.8,1557.5,2109.2,1269.4,2543.9,472.45,1689.7,358.41,642.71,739.26,0.0000,-3533.8,-6576.2,-293.71,-2708.6,-2498.0,-13691.,-1684.2,-1300.0,-5186.8,-2786.4,-5704.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1319.000000000,6361.8,1435.7,1544.8,1563.1,2099.9,1277.5,2493.0,474.83,1694.5,358.92,643.80,748.54,0.0000,-3530.2,-6573.2,-293.30,-2707.5,-2496.5,-13688.,-1684.1,-1298.5,-5186.2,-2785.8,-5703.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1320.000000000,6347.2,1453.0,1546.6,1573.4,2110.6,1234.1,2509.9,474.74,1679.5,363.02,642.60,755.80,0.0000,-3526.7,-6570.1,-292.91,-2706.4,-2495.0,-13686.,-1684.1,-1297.1,-5185.1,-2785.2,-5702.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1321.000000000,6389.3,1440.4,1531.2,1574.7,2119.1,1215.1,2474.1,476.76,1688.5,368.76,640.75,762.11,0.0000,-3566.7,-6588.4,-296.53,-2705.4,-2521.2,-13685.,-1704.5,-1313.9,-5200.0,-2787.2,-5715.0,0.15344E+06,68585.,52538.,49309.,95587.,32939.,0.11807E+06,34119.,52159.,15569.,22375.,26952.,0.0000,-154.94,-161.32,-24.841,-148.04,-96.179,-601.21,-485.74,-49.681,-436.36,-52.804,-592.44
1322.000000000,6406.0,1439.0,1511.6,1576.5,2100.8,1211.7,2459.4,480.32,1716.3,365.53,630.14,760.73,0.0000,-3585.8,-6609.3,-300.00,-2704.6,-2530.6,-13683.,-1717.2,-1325.9,-5208.7,-2787.8,-5724.5,0.13271E+06,59320.,45440.,42647.,82674.,28489.,0.10212E+06,29509.,45113.,13466.,19352.,23311.,0.0000,-134.24,-139.61,-21.485,-128.13,-83.298,-519.98,-420.20,-42.970,-377.41,-45.672,-512.40
1323.000000000,6538.9,1430.5,1543.1,1586.5,2102.4,1224.0,2511.7,479.37,1747.8,369.58,630.62,776.78,0.0000,-3601.3,-6628.8,-302.77,-2704.2,-2538.5,-13683.,-1715.2,-1335.6,-5212.9,-2788.3,-5729.3,50635.,22633.,17337.,16272.,31543.,10870.,38962.,11259.,17212.,5137.7,7383.8,8894.1,0.0000,-51.332,-53.324,-8.1973,-48.944,-31.858,-198.49,-160.37,-16.395,-144.01,-17.427,-195.57
1324.000000000,6560.7,1494.0,1587.1,1594.2,2128.2,1294.2,2524.7,486.68,1780.6,375.86,650.61,786.16,0.0000,-3619.5,-6649.9,-304.97,-2704.8,-2547.9,-13687.,-1708.1,-1343.8,-5214.2,-2790.3,-5730.1,10191.,4555.0,3489.3,3274.8,6348.3,2187.6,7841.3,2266.0,3464.1,1034.0,1486.0,1790.0,0.0000,-10.378,-10.746,-1.6498,-9.8723,-6.4444,-39.987,-32.290,-3.2995,-28.992,-3.5102,-39.385
1325.000000000,6578.6,1451.8,1657.2,1587.8,2113.2,1261.7,2460.8,468.92,1797.7,375.39,643.73,790.08,0.0000,-3634.2,-6668.6,-306.73,-2704.7,-2554.0,-13690.,-1713.8,-1351.1,-5217.2,-2791.0,-5732.0,93503.,41794.,32015.,30047.,58248.,20072.,71947.,20791.,31784.,9487.3,13635.,16424.,0.0000,-95.448,-98.686,-15.137,-90.692,-59.240,-366.98,-296.37,-30.275,-266.05,-32.208,-361.50
1326.000000000,6542.2,1446.7,1672.6,1603.2,2135.1,1242.7,2443.1,464.37,1813.8,366.70,644.86,792.47,0.0000,-3647.9,-6684.2,-308.18,-2705.1,-2559.3,-13693.,-1709.5,-1357.9,-5218.1,-2792.2,-5732.5,28843.,12892.,9875.7,9268.7,17968.,6191.6,22194.,6413.4,9804.5,2926.5,4205.9,5066.3,0.0000,-29.508,-30.467,-4.6694,-28.001,-18.296,-113.21,-91.443,-9.3387,-82.078,-9.9358,-111.54
1327.000000000,6542.6,1480.1,1673.8,1594.9,2187.3,1295.9,2461.8,476.29,1847.4,366.32,647.19,801.83,0.0000,-3661.3,-6697.7,-309.42,-2705.8,-2565.3,-13695.,-1704.0,-1364.3,-5217.4,-2793.3,-5731.6,11133.,4976.2,3811.9,3577.6,6935.3,2389.9,8566.3,2475.5,3784.4,1129.6,1623.4,1955.5,0.0000,-11.419,-11.772,-1.8023,-10.820,-7.0767,-43.713,-35.305,-3.6046,-31.686,-3.8357,-43.072
1328.000000000,6619.5,1471.7,1670.2,1572.9,2180.9,1281.9,2470.6,466.96,1850.6,366.16,650.24,806.14,0.0000,-3673.9,-6710.4,-310.53,-2706.0,-2570.5,-13699.,-1741.7,-1370.2,-5225.6,-2794.5,-5741.4,0.32257E+06,0.14418E+06,0.11045E+06,0.10366E+06,0.20094E+06,69244.,0.24820E+06,71725.,0.10965E+06,32729.,47038.,56659.,0.0000,-331.59,-341.38,-52.220,-313.75,-205.23,-1266.7,-1023.5,-104.44,-918.21,-111.15,-1248.4
1329.000000000,6730.1,1651.4,1746.0,1563.7,2271.2,1415.3,2657.5,487.68,1778.1,399.34,716.15,884.01,0.0000,-3694.0,-6729.5,-311.82,-2708.9,-2583.5,-13710.,-1732.2,-1376.0,-5234.1,-2801.5,-5746.5,40588.,18142.,13897.,13043.,25284.,8712.9,31231.,9025.0,13797.,4118.3,5918.7,7129.3,0.0000,-42.009,-43.056,-6.5708,-39.624,-26.097,-159.80,-128.94,-13.142,-115.63,-14.010,-157.38
1330.000000000,6749.2,1723.4,1747.2,1554.6,2317.2,1294.3,2548.1,499.56,1791.9,406.33,781.45,908.58,0.0000,-3711.2,-6744.1,-313.21,-2712.0,-2589.5,-13717.,-1727.6,-1381.9,-5240.3,-2813.7,-5749.1,62330.,27860.,21342.,20030.,38829.,13380.,47961.,13859.,21188.,6324.3,9089.1,10948.,0.0000,-64.657,-66.165,-10.091,-60.906,-40.131,-245.41,-198.10,-20.181,-177.61,-21.526,-241.82
1331.000000000,6821.0,1739.4,1713.6,1562.0,2399.4,1266.3,2548.2,524.50,1815.3,391.21,825.82,885.98,0.0000,-3724.1,-6759.0,-314.60,-2711.6,-2593.5,-13721.,-1725.9,-1387.6,-5240.5,-2824.9,-5751.2,76361.,34132.,26146.,24539.,47569.,16392.,58757.,16979.,25957.,7747.9,11135.,13413.,0.0000,-79.294,-81.104,-12.362,-74.636,-49.106,-300.54,-242.76,-24.724,-217.61,-26.376,-296.32
1332.000000000,6778.4,1718.1,1662.9,1553.9,2426.5,1226.2,2672.1,535.19,1770.9,387.38,758.51,856.84,0.0000,-3692.9,-6742.3,-311.85,-2710.3,-2569.9,-13723.,-1714.5,-1368.2,-5225.3,-2824.6,-5741.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1333.000000000,6823.1,1741.5,1655.2,1591.2,2423.4,1261.1,2744.8,535.10,1750.2,406.54,731.03,846.73,0.0000,-3728.1,-6746.9,-313.24,-2709.3,-2591.3,-13728.,-1707.5,-1381.8,-5231.4,-2825.4,-5744.3,10090.,4509.9,3454.7,3242.4,6285.5,2165.9,7763.7,2243.5,3429.8,1023.8,1471.3,1772.3,0.0000,-10.492,-10.728,-1.6334,-9.8639,-6.4862,-39.722,-32.093,-3.2669,-28.762,-3.4859,-39.182
1334.000000000,6651.1,1790.0,1655.7,1587.1,2403.2,1242.9,2710.3,512.36,1725.4,412.83,702.75,861.43,0.0000,-3700.0,-6732.3,-310.94,-2708.7,-2568.6,-13729.,-1701.2,-1365.0,-5219.7,-2821.5,-5735.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1335.000000000,6561.0,1761.0,1700.5,1603.1,2516.0,1215.0,2659.1,511.78,1725.5,414.05,700.66,859.11,0.0000,-3688.7,-6716.3,-308.67,-2707.9,-2561.1,-13730.,-1696.7,-1356.1,-5214.5,-2819.5,-5731.7,37.258,16.654,12.757,11.973,23.210,7.9981,28.669,8.2846,12.665,3.7804,5.4331,6.5445,0.0000,-0.38658E-01,-0.39605E-01,-0.60318E-02,-0.36360E-01,-0.23838E-01,-0.14659,-0.11852,-0.12064E-01,-0.10622,-0.12865E-01,-0.14470
1336.000000000,6531.4,1751.1,1734.5,1607.9,2523.2,1215.9,2592.9,502.33,1709.3,405.90,721.43,860.61,0.0000,-3724.5,-6725.6,-310.92,-2707.2,-2584.0,-13731.,-1694.3,-1372.8,-5222.5,-2823.1,-5737.6,5242.8,2343.4,1795.1,1684.8,3266.0,1125.5,4034.2,1165.8,1782.2,531.96,764.52,920.91,0.0000,-5.4455,-5.5752,-0.84876,-5.1193,-3.3569,-20.620,-16.677,-1.6975,-14.947,-1.8099,-20.361
1337.000000000,6576.3,1717.2,1735.8,1580.8,2469.8,1238.0,2663.8,501.73,1728.3,405.98,707.24,860.21,0.0000,-3740.0,-6738.5,-313.39,-2707.2,-2590.9,-13732.,-1695.1,-1382.2,-5224.8,-2824.6,-5740.1,23293.,10412.,7975.6,7485.4,14511.,5000.3,17923.,5179.4,7918.1,2363.5,3396.7,4091.5,0.0000,-24.232,-24.789,-3.7710,-22.763,-14.924,-91.599,-74.093,-7.5420,-66.407,-8.0400,-90.456
1338.000000000,6592.1,1678.1,1743.9,1572.5,2424.0,1251.1,2656.4,496.79,1748.4,400.25,693.64,854.54,0.0000,-3753.7,-6751.5,-315.42,-2707.1,-2595.5,-13734.,-1694.1,-1390.4,-5225.7,-2823.5,-5741.1,10359.,4630.2,3546.8,3328.8,6453.1,2223.7,7970.8,2303.4,3521.3,1051.1,1510.6,1819.5,0.0000,-10.795,-11.033,-1.6770,-10.130,-6.6385,-40.729,-32.948,-3.3540,-29.531,-3.5750,-40.222
1339.000000000,6566.9,1642.2,1757.7,1555.3,2463.9,1265.0,2645.5,489.76,1742.2,395.60,694.04,830.18,0.0000,-3765.7,-6762.3,-317.03,-2707.6,-2599.7,-13736.,-1695.0,-1396.5,-5227.2,-2821.8,-5741.8,21873.,9777.0,7489.4,7029.1,13626.,4695.5,16831.,4863.7,7435.4,2219.4,3189.6,3842.1,0.0000,-22.830,-23.317,-3.5411,-21.403,-14.020,-85.987,-69.567,-7.0822,-62.355,-7.5474,-84.921
1340.000000000,6503.8,1619.7,1710.1,1548.3,2498.3,1302.7,2646.0,478.59,1796.2,403.81,691.16,825.78,0.0000,-3775.9,-6771.9,-318.32,-2709.6,-2604.1,-13736.,-1694.4,-1401.5,-5227.8,-2821.0,-5742.5,12926.,5777.8,4426.0,4153.9,8052.5,2774.9,9946.4,2874.3,4394.0,1311.6,1885.0,2270.5,0.0000,-13.514,-13.792,-2.0926,-12.656,-8.2884,-50.811,-41.109,-4.1853,-36.848,-4.4595,-50.179
1341.000000000,6561.1,1622.6,1681.4,1591.8,2487.2,1346.2,2700.9,474.33,1788.5,404.24,678.64,825.35,0.0000,-3786.7,-6781.9,-319.39,-2711.2,-2608.3,-13736.,-1693.9,-1406.4,-5227.4,-2819.6,-5742.9,12928.,5778.8,4426.7,4154.6,8053.9,2775.3,9948.0,2874.7,4394.8,1311.8,1885.3,2270.9,0.0000,-13.540,-13.806,-2.0930,-12.666,-8.2941,-50.817,-41.113,-4.1860,-36.853,-4.4597,-50.181
1342.000000000,6519.6,1633.9,1660.8,1618.6,2544.2,1316.1,2700.6,471.43,1828.8,410.44,668.59,814.61,0.0000,-3796.9,-6791.1,-320.32,-2713.6,-2612.6,-13736.,-1698.1,-1410.6,-5228.9,-2818.2,-5743.8,46384.,20733.,15882.,14906.,28895.,9957.2,35691.,10314.,15767.,4706.4,6763.9,8147.5,0.0000,-48.663,-49.577,-7.5092,-45.470,-29.775,-182.32,-147.50,-15.018,-132.21,-15.999,-180.02
1343.000000000,6542.4,1648.0,1681.2,1621.5,2564.1,1326.8,2631.2,474.16,1859.0,412.66,675.11,808.83,0.0000,-3760.7,-6776.7,-317.09,-2715.9,-2589.6,-13735.,-1695.0,-1389.2,-5217.5,-2814.2,-5735.4,772.00,345.07,264.33,248.08,480.92,165.72,594.03,171.66,262.43,78.331,112.58,135.60,0.0000,-0.80933,-0.82531,-0.12498,-0.75600,-0.49462,-3.0345,-2.4547,-0.24996,-2.2004,-0.26623,-2.9958
1344.000000000,6489.9,1638.8,1684.4,1619.8,2583.2,1320.4,2545.4,470.60,1890.6,412.23,692.41,810.75,0.0000,-3745.9,-6759.1,-314.00,-2718.1,-2583.6,-13735.,-1692.5,-1377.5,-5213.3,-2812.6,-5731.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1345.000000000,6663.5,1659.4,1712.7,1605.2,2571.6,1332.4,2546.6,471.06,1876.7,407.85,701.07,817.13,0.0000,-3735.0,-6742.6,-311.61,-2719.8,-2579.9,-13735.,-1690.7,-1369.0,-5209.8,-2812.0,-5728.4,367.31,164.18,125.77,118.04,228.82,78.849,282.63,81.673,124.86,37.269,53.562,64.518,0.0000,-0.38434,-0.39258,-0.59464E-01,-0.35934,-0.23516,-1.4442,-1.1679,-0.11893,-1.0469,-0.12666,-1.4253
1346.000000000,6676.7,1655.1,1697.2,1594.9,2580.4,1336.6,2578.4,464.33,1853.9,404.87,703.50,809.57,0.0000,-3725.7,-6728.0,-309.79,-2721.0,-2576.7,-13737.,-1689.4,-1362.3,-5207.6,-2811.5,-5726.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1347.000000000,6693.3,1679.2,1689.5,1577.3,2546.3,1323.6,2591.3,451.04,1791.7,397.86,695.61,818.59,0.0000,-3716.7,-6713.9,-308.36,-2721.4,-2572.9,-13737.,-1688.4,-1356.6,-5206.5,-2810.8,-5724.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1348.000000000,6615.5,1629.0,1672.5,1589.9,2549.0,1323.1,2639.9,445.67,1805.4,391.20,691.89,807.99,0.0000,-3708.5,-6701.2,-307.21,-2722.0,-2569.1,-13739.,-1687.7,-1351.6,-5205.6,-2809.3,-5723.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1349.000000000,6585.6,1585.2,1651.0,1603.8,2506.0,1315.6,2612.0,452.81,1830.5,388.87,694.22,792.53,0.0000,-3700.9,-6690.5,-306.26,-2722.8,-2565.4,-13739.,-1687.2,-1347.3,-5204.4,-2807.8,-5722.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1350.000000000,6578.6,1584.2,1673.6,1618.0,2484.8,1331.8,2648.8,457.10,1815.7,387.36,700.53,779.75,0.0000,-3738.6,-6706.1,-309.48,-2723.6,-2590.2,-13740.,-1689.1,-1365.3,-5215.3,-2808.8,-5729.3,16292.,7282.4,5578.5,5235.6,10149.,3497.5,12537.,3622.7,5538.3,1653.1,2375.8,2861.8,0.0000,-16.991,-17.389,-2.6376,-15.933,-10.431,-64.064,-51.789,-5.2752,-46.430,-5.6173,-63.197
1351.000000000,6654.4,1581.8,1672.7,1608.8,2515.4,1332.7,2650.8,456.30,1758.6,379.44,705.42,782.26,0.0000,-3709.6,-6700.1,-308.58,-2724.3,-2570.3,-13740.,-1688.3,-1353.1,-5206.7,-2806.5,-5723.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1352.000000000,6658.2,1587.7,1656.1,1616.9,2489.6,1335.9,2641.0,463.61,1746.5,382.70,702.65,790.40,0.0000,-3744.0,-6714.0,-311.31,-2724.5,-2592.9,-13742.,-1693.4,-1369.2,-5216.5,-2808.0,-5730.9,42130.,18832.,14425.,13539.,26245.,9044.0,32418.,9368.0,14321.,4274.8,6143.6,7400.3,0.0000,-43.958,-44.976,-6.8205,-41.229,-26.981,-165.63,-133.90,-13.641,-120.05,-14.527,-163.38
1353.000000000,6797.9,1581.6,1605.3,1634.2,2448.1,1323.6,2633.3,463.20,1779.7,383.17,695.87,781.39,0.0000,-3758.8,-6729.2,-314.02,-2724.8,-2600.2,-13742.,-1692.1,-1379.1,-5219.4,-2808.4,-5733.2,3910.8,1748.1,1339.1,1256.8,2436.3,839.53,3009.3,869.61,1329.4,396.81,570.29,686.95,0.0000,-4.0865,-4.1773,-0.63313,-3.8308,-2.5069,-15.373,-12.429,-1.2663,-11.144,-1.3486,-15.164
1354.000000000,6825.5,1607.7,1586.3,1639.6,2409.0,1301.7,2661.0,468.92,1805.1,386.13,689.25,800.13,0.0000,-3770.2,-6742.9,-316.22,-2725.0,-2605.7,-13741.,-1693.0,-1386.7,-5220.8,-2809.0,-5734.4,18706.,8361.4,6405.1,6011.4,11653.,4015.7,14394.,4159.5,6358.9,1898.0,2727.8,3285.8,0.0000,-19.577,-19.994,-3.0284,-18.339,-12.000,-73.523,-59.445,-6.0568,-53.302,-6.4509,-72.525
1355.000000000,6827.7,1574.8,1576.7,1640.6,2262.6,1246.1,2657.4,468.74,1788.8,377.90,694.34,803.79,0.0000,-3734.9,-6731.9,-313.90,-2724.7,-2582.2,-13739.,-1691.1,-1369.1,-5209.7,-2806.7,-5726.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1356.000000000,6837.2,1567.8,1588.3,1661.2,2260.1,1255.6,2654.1,462.85,1765.0,376.53,684.81,787.27,0.0000,-3720.9,-6717.6,-311.45,-2724.2,-2575.4,-13738.,-1689.6,-1360.2,-5205.5,-2805.2,-5723.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1357.000000000,6894.8,1584.7,1585.4,1689.7,2236.3,1275.3,2648.6,461.40,1803.3,379.51,681.34,777.41,0.0000,-3710.2,-6704.4,-309.47,-2723.7,-2570.8,-13737.,-1688.5,-1353.7,-5203.2,-2804.0,-5722.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1358.000000000,6918.5,1589.1,1575.5,1669.7,2219.9,1250.1,2705.2,466.42,1811.6,371.70,674.58,778.89,0.0000,-3700.8,-6692.2,-307.93,-2723.2,-2566.8,-13738.,-1687.6,-1348.4,-5201.7,-2802.8,-5720.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1359.000000000,6954.3,1589.8,1589.6,1641.0,2229.0,1251.5,2701.4,474.73,1796.9,370.49,662.77,777.00,0.0000,-3692.3,-6681.5,-306.72,-2722.7,-2563.4,-13738.,-1687.1,-1343.9,-5200.5,-2801.8,-5719.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1360.000000000,6984.6,1593.0,1626.1,1630.6,2225.7,1290.7,2748.2,471.78,1784.8,369.18,654.05,769.67,0.0000,-3684.6,-6672.3,-305.75,-2722.1,-2560.2,-13739.,-1686.6,-1340.2,-5199.6,-2801.1,-5718.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1361.000000000,6909.5,1593.4,1586.6,1645.4,2312.2,1278.6,2750.6,468.95,1772.3,373.79,651.16,767.32,0.0000,-3677.5,-6663.1,-304.93,-2721.4,-2557.1,-13739.,-1686.3,-1336.9,-5198.9,-2800.5,-5717.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1362.000000000,6907.8,1609.9,1594.1,1628.1,2275.0,1276.6,2733.5,465.80,1785.5,370.81,641.39,764.62,0.0000,-3670.8,-6655.3,-304.23,-2720.6,-2553.9,-13739.,-1686.1,-1333.9,-5198.3,-2799.6,-5717.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1363.000000000,6720.8,1620.6,1622.7,1627.7,2231.9,1285.0,2725.3,466.99,1797.2,366.44,641.98,761.08,0.0000,-3664.4,-6648.2,-303.60,-2719.8,-2550.8,-13739.,-1685.9,-1331.2,-5197.6,-2798.8,-5716.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1364.000000000,6596.1,1641.1,1627.5,1620.8,2208.9,1317.3,2671.2,464.17,1791.4,365.40,636.45,764.65,0.0000,-3703.1,-6664.8,-307.04,-2719.2,-2575.8,-13739.,-1712.9,-1349.8,-5213.8,-2800.4,-5731.0,0.20247E+06,90501.,69326.,65065.,0.12613E+06,43464.,0.15580E+06,45021.,68826.,20544.,29525.,35564.,0.0000,-209.99,-215.75,-32.778,-197.68,-129.07,-795.38,-643.04,-65.557,-576.71,-69.793,-784.12
1365.000000000,6787.9,1700.9,1626.7,1609.8,2215.1,1387.1,2801.8,475.21,1797.8,379.86,635.30,785.68,0.0000,-3722.0,-6683.3,-310.39,-2720.0,-2587.4,-13741.,-1769.0,-1361.6,-5232.9,-2801.6,-5753.7,0.46535E+06,0.20800E+06,0.15934E+06,0.14954E+06,0.28989E+06,99896.,0.35807E+06,0.10347E+06,0.15819E+06,47217.,67859.,81740.,0.0000,-484.17,-496.49,-75.336,-455.37,-298.23,-1830.5,-1479.5,-150.67,-1325.9,-160.46,-1803.9
1366.000000000,6805.3,2109.5,1843.6,1622.6,2359.0,1630.4,3110.9,487.55,1798.3,457.75,799.12,918.04,0.0000,-3756.4,-6717.5,-313.31,-2727.5,-2607.3,-13760.,-1754.2,-1370.8,-5254.3,-2816.0,-5765.4,50996.,22794.,17461.,16388.,31768.,10947.,39240.,11339.,17335.,5174.3,7436.4,8957.5,0.0000,-53.632,-54.562,-8.2557,-50.193,-33.269,-201.44,-162.41,-16.511,-145.47,-17.644,-198.21
1367.000000000,6824.7,2064.5,1742.9,1627.6,2346.7,1397.6,2847.2,493.86,1841.1,423.01,836.43,904.62,0.0000,-3730.2,-6715.4,-311.78,-2731.0,-2584.8,-13765.,-1735.6,-1356.3,-5247.0,-2826.7,-5759.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1368.000000000,6732.7,2078.3,1726.9,1658.4,2366.3,1359.3,2818.4,508.16,1846.7,407.16,861.67,870.87,0.0000,-3720.6,-6709.1,-310.04,-2730.7,-2577.8,-13768.,-1721.4,-1350.0,-5239.3,-2836.3,-5754.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1369.000000000,6713.7,2021.5,1701.6,1691.9,2344.7,1354.1,2991.3,536.99,1835.8,408.36,796.71,838.85,0.0000,-3715.7,-6697.3,-308.67,-2729.2,-2572.4,-13770.,-1711.2,-1345.8,-5232.5,-2836.9,-5748.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1370.000000000,6654.9,2020.7,1682.1,1699.4,2344.4,1364.0,3016.5,518.63,1802.1,413.71,748.37,832.49,0.0000,-3711.3,-6685.5,-307.60,-2727.6,-2567.3,-13772.,-1704.0,-1342.4,-5228.0,-2833.6,-5744.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1371.000000000,6654.3,1954.7,1777.4,1680.4,2419.8,1357.2,2966.2,505.84,1819.6,419.62,730.47,837.76,0.0000,-3705.9,-6675.8,-306.74,-2726.7,-2562.7,-13773.,-1699.0,-1339.5,-5224.8,-2829.7,-5742.1,9.0637,4.0513,3.1034,2.9126,5.6463,1.9457,6.9742,2.0154,3.0810,0.91965,1.3217,1.5920,0.0000,-0.94516E-02,-0.96751E-02,-0.14673E-02,-0.88773E-02,-0.58467E-02,-0.35728E-01,-0.28883E-01,-0.29346E-02,-0.25863E-01,-0.31330E-02,-0.35255E-01
1372.000000000,6560.6,1902.6,1788.4,1657.7,2441.5,1383.4,2916.5,497.08,1786.5,409.62,756.13,848.52,0.0000,-3699.1,-6668.6,-306.02,-2726.2,-2558.9,-13773.,-1695.6,-1336.7,-5222.3,-2829.7,-5740.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1373.000000000,6587.5,1843.6,1799.0,1636.6,2357.6,1377.2,2939.1,498.25,1801.5,409.42,746.49,851.20,0.0000,-3692.6,-6665.1,-305.39,-2726.1,-2555.8,-13772.,-1693.3,-1335.5,-5221.4,-2829.7,-5739.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1374.000000000,6700.1,1839.9,1818.6,1623.0,2399.6,1348.0,2952.4,490.41,1782.7,407.00,737.62,842.08,0.0000,-3688.7,-6659.7,-304.82,-2726.8,-2553.3,-13773.,-1691.7,-1334.4,-5221.5,-2827.7,-5737.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1375.000000000,6688.4,1866.3,1771.3,1616.4,2465.5,1399.5,2918.8,484.94,1805.5,411.74,737.06,822.41,0.0000,-3684.1,-6654.9,-304.28,-2728.4,-2551.0,-13773.,-1690.5,-1332.3,-5221.0,-2825.5,-5735.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1376.000000000,6661.6,1828.4,1793.9,1612.7,2408.1,1394.7,2920.8,484.95,1747.8,404.00,721.77,806.95,0.0000,-3679.8,-6653.4,-303.77,-2729.2,-2548.7,-13772.,-1689.7,-1330.3,-5219.4,-2823.4,-5734.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1377.000000000,6633.5,1794.0,1773.1,1584.5,2411.5,1431.9,2926.1,476.80,1749.6,403.85,721.54,807.56,0.0000,-3675.1,-6650.1,-303.28,-2730.7,-2547.4,-13771.,-1689.3,-1328.5,-5218.3,-2822.1,-5733.2,1016.3,454.27,347.98,326.59,633.12,218.17,782.02,225.98,345.47,103.12,148.20,178.52,0.0000,-1.0532,-1.0833,-0.16453,-0.99264,-0.65214,-4.0028,-3.2367,-0.32906,-2.8992,-0.35080,-3.9496
1378.000000000,6617.4,1803.8,1748.8,1565.0,2388.4,1439.6,2886.4,475.22,1770.2,405.44,719.56,806.13,0.0000,-3670.8,-6646.2,-302.80,-2732.2,-2546.0,-13770.,-1688.8,-1326.8,-5217.2,-2821.0,-5732.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1379.000000000,6419.5,1800.3,1752.3,1555.2,2400.7,1419.5,2849.0,469.67,1749.0,409.36,734.73,796.73,0.0000,-3666.4,-6641.9,-302.34,-2733.4,-2544.4,-13768.,-1688.5,-1325.0,-5215.9,-2819.9,-5731.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1380.000000000,6417.2,1800.9,1725.1,1573.8,2387.3,1402.4,2852.4,469.43,1737.8,406.90,741.73,790.42,0.0000,-3661.9,-6637.2,-301.90,-2734.5,-2542.7,-13768.,-1688.2,-1323.3,-5214.4,-2818.9,-5730.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1381.000000000,6421.4,1810.0,1713.8,1577.1,2354.8,1393.5,2822.3,473.73,1760.9,406.75,736.14,792.86,0.0000,-3657.4,-6632.3,-301.48,-2735.1,-2541.0,-13768.,-1688.0,-1321.9,-5213.2,-2817.8,-5729.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1382.000000000,6507.0,1778.2,1688.7,1569.9,2323.9,1389.8,2813.3,475.93,1791.1,405.23,740.07,789.15,0.0000,-3652.7,-6627.1,-301.06,-2735.5,-2539.2,-13767.,-1687.9,-1320.7,-5212.1,-2816.6,-5728.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1383.000000000,6686.7,1778.1,1712.8,1571.9,2323.0,1391.4,2815.2,475.54,1813.0,407.05,748.33,789.43,0.0000,-3648.0,-6624.4,-300.66,-2735.8,-2537.0,-13767.,-1687.7,-1319.3,-5211.5,-2815.5,-5727.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1384.000000000,6674.0,1765.0,1748.4,1567.0,2322.6,1405.3,2767.2,476.03,1802.3,407.76,755.59,794.50,0.0000,-3643.3,-6623.3,-300.27,-2736.0,-2535.1,-13767.,-1687.6,-1318.1,-5210.8,-2814.7,-5727.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1385.000000000,6597.4,1753.9,1762.8,1563.7,2320.8,1368.9,2741.6,469.14,1807.7,408.92,748.20,801.53,0.0000,-3638.6,-6621.8,-299.88,-2736.0,-2533.1,-13768.,-1687.5,-1317.0,-5210.3,-2814.0,-5727.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1386.000000000,6590.8,1730.2,1753.1,1560.6,2323.7,1370.7,2732.1,465.92,1823.4,407.07,753.22,798.18,0.0000,-3633.9,-6619.5,-299.52,-2736.0,-2531.3,-13768.,-1687.5,-1316.1,-5210.0,-2813.3,-5726.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1387.000000000,6611.3,1717.7,1772.6,1562.7,2305.0,1382.1,2739.8,469.65,1862.4,401.34,756.05,808.04,0.0000,-3629.3,-6616.2,-299.16,-2735.7,-2529.4,-13767.,-1687.4,-1315.1,-5209.7,-2812.7,-5726.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1388.000000000,6649.3,1713.4,1766.3,1585.3,2292.7,1359.8,2734.1,468.28,1882.2,396.98,740.88,809.88,0.0000,-3624.9,-6613.1,-298.84,-2735.2,-2527.5,-13768.,-1687.3,-1314.1,-5209.3,-2811.6,-5726.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1389.000000000,6739.6,1708.7,1746.7,1596.8,2293.7,1353.0,2722.0,469.32,1878.6,398.20,730.75,808.56,0.0000,-3620.6,-6610.4,-298.56,-2734.7,-2525.7,-13768.,-1687.3,-1313.2,-5208.7,-2810.4,-5726.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1390.000000000,6999.7,1732.9,1718.0,1578.8,2318.9,1351.8,2728.8,461.75,1854.4,402.99,731.86,800.94,0.0000,-3616.3,-6607.2,-298.29,-2734.1,-2523.8,-13770.,-1687.3,-1312.3,-5208.0,-2809.1,-5725.8,856.54,382.86,293.28,275.25,533.59,183.87,659.08,190.46,291.16,86.909,124.90,150.45,0.0000,-0.87785,-0.90902,-0.13867,-0.83367,-0.54657,-3.3714,-2.7238,-0.27733,-2.4415,-0.29549,-3.3214
1391.000000000,7060.9,1732.1,1816.4,1599.6,2289.1,1364.7,2761.2,464.52,1859.5,409.86,725.26,791.93,0.0000,-3612.2,-6603.8,-298.02,-2733.5,-2521.9,-13770.,-1687.2,-1311.5,-5207.3,-2808.1,-5725.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1392.000000000,7093.0,1737.2,1832.8,1603.7,2267.5,1373.6,2783.4,462.84,1836.8,406.82,716.17,786.65,0.0000,-3607.9,-6601.0,-297.75,-2732.9,-2520.2,-13770.,-1687.2,-1310.7,-5206.7,-2807.2,-5725.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1393.000000000,6947.5,1764.9,1844.1,1598.2,2249.0,1372.7,2798.3,456.71,1844.2,405.51,709.83,787.03,0.0000,-3603.7,-6597.4,-297.48,-2732.0,-2518.4,-13768.,-1687.1,-1309.9,-5205.8,-2806.4,-5724.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1394.000000000,6836.2,1788.1,1859.4,1613.5,2217.7,1369.8,2783.7,455.37,1839.0,407.08,701.03,791.87,0.0000,-3599.5,-6594.3,-297.19,-2731.0,-2516.6,-13767.,-1687.1,-1309.0,-5205.1,-2805.7,-5724.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1395.000000000,6862.1,1774.6,1861.0,1638.4,2232.4,1371.8,2768.6,454.46,1840.5,404.13,696.74,791.91,0.0000,-3595.3,-6591.4,-296.88,-2729.9,-2514.8,-13765.,-1687.0,-1308.1,-5204.4,-2805.1,-5724.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1396.000000000,6904.2,1780.7,1848.7,1619.5,2234.7,1366.1,2785.3,453.37,1844.2,402.14,694.61,784.41,0.0000,-3591.1,-6588.3,-296.55,-2729.6,-2513.1,-13764.,-1686.9,-1307.5,-5204.1,-2804.5,-5724.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1397.000000000,7110.0,1819.3,1809.9,1637.6,2206.2,1362.7,2764.5,453.22,1846.1,397.23,702.57,773.59,0.0000,-3587.0,-6585.5,-296.26,-2728.9,-2511.4,-13763.,-1686.9,-1306.9,-5203.7,-2804.0,-5723.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1398.000000000,7215.4,1808.5,1814.6,1623.8,2187.9,1371.8,2792.2,451.20,1849.9,392.66,710.79,770.95,0.0000,-3583.0,-6583.0,-295.97,-2728.1,-2509.5,-13761.,-1686.8,-1306.3,-5203.4,-2803.3,-5723.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1399.000000000,7166.3,1778.5,1802.0,1595.4,2197.9,1375.2,2770.9,452.66,1841.1,384.45,721.76,771.19,0.0000,-3579.1,-6580.8,-295.68,-2727.3,-2507.8,-13759.,-1686.8,-1305.8,-5202.9,-2802.6,-5722.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1400.000000000,7084.9,1739.1,1798.9,1608.4,2110.9,1384.6,2768.1,448.77,1855.0,383.17,722.94,768.24,0.0000,-3575.3,-6579.6,-295.38,-2726.5,-2506.1,-13756.,-1686.7,-1305.2,-5202.8,-2801.9,-5722.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1401.000000000,6993.1,1736.0,1785.7,1623.7,2008.8,1415.8,2779.3,451.24,1834.8,386.64,727.54,769.14,0.0000,-3571.5,-6578.6,-295.09,-2725.7,-2504.5,-13754.,-1686.7,-1304.6,-5202.6,-2801.2,-5722.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1402.000000000,6807.3,1742.4,1808.4,1622.4,2000.5,1408.8,2761.4,460.66,1846.2,391.47,725.88,774.36,0.0000,-3567.8,-6577.3,-294.79,-2724.9,-2503.0,-13751.,-1686.6,-1303.9,-5202.4,-2800.6,-5721.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1403.000000000,6817.9,1739.4,1828.5,1631.6,2024.5,1421.3,2759.3,460.09,1846.6,390.95,720.55,778.42,0.0000,-3564.3,-6576.0,-294.49,-2724.0,-2501.7,-13748.,-1686.5,-1303.2,-5202.1,-2800.1,-5721.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1404.000000000,6792.6,1759.1,1863.6,1667.9,2093.0,1443.2,2789.8,455.94,1881.0,389.55,727.17,776.36,0.0000,-3604.8,-6597.9,-298.19,-2723.2,-2528.2,-13747.,-1698.4,-1320.9,-5215.8,-2802.3,-5731.4,88814.,39698.,30410.,28541.,55327.,19066.,68340.,19749.,30191.,9011.6,12951.,15600.,0.0000,-90.301,-93.848,-14.378,-86.064,-56.287,-349.28,-282.01,-28.756,-252.96,-30.622,-343.60
1405.000000000,6710.8,1811.0,1864.0,1654.3,2097.9,1458.1,2782.1,459.41,1909.3,391.55,734.40,780.75,0.0000,-3624.2,-6621.5,-301.72,-2722.5,-2538.0,-13745.,-1695.9,-1333.8,-5220.4,-2803.0,-5734.9,3167.1,1415.6,1084.4,1017.7,1972.9,679.87,2437.0,704.22,1076.6,321.35,461.83,556.30,0.0000,-3.2271,-3.3487,-0.51272,-3.0710,-2.0096,-12.455,-10.056,-1.0254,-9.0199,-1.0920,-12.251
1406.000000000,6630.8,1832.4,1849.3,1651.3,2065.9,1442.6,2759.6,458.20,1918.6,396.75,732.36,784.56,0.0000,-3640.1,-6642.6,-304.56,-2721.6,-2545.4,-13743.,-1693.6,-1344.1,-5221.5,-2803.4,-5735.6,1506.0,673.16,515.65,483.96,938.18,323.29,1158.8,334.87,511.94,152.81,219.61,264.53,0.0000,-1.5380,-1.5936,-0.24381,-1.4618,-0.95641,-5.9223,-4.7814,-0.48762,-4.2890,-0.51929,-5.8249
1407.000000000,6576.4,1806.3,1846.2,1649.1,2060.5,1425.8,2771.4,456.37,1906.5,396.43,719.49,785.95,0.0000,-3654.4,-6661.5,-306.79,-2720.8,-2552.0,-13741.,-1693.2,-1353.0,-5221.6,-2803.4,-5735.5,11887.,5313.1,4070.0,3819.8,7404.9,2551.7,9146.4,2643.1,4040.6,1206.1,1733.4,2087.9,0.0000,-12.166,-12.588,-1.9243,-11.548,-7.5537,-46.743,-37.736,-3.8487,-33.851,-4.0987,-45.970
1408.000000000,6609.9,1790.3,1828.7,1618.3,2015.4,1417.3,2785.0,457.30,1907.1,397.51,712.45,779.90,0.0000,-3622.9,-6655.0,-304.55,-2719.7,-2530.2,-13739.,-1691.3,-1338.8,-5209.7,-2800.6,-5726.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1409.000000000,6742.3,1744.2,1831.5,1603.5,2034.4,1400.4,2805.7,460.11,1932.4,395.13,705.79,769.88,0.0000,-3612.0,-6645.0,-302.19,-2718.5,-2524.8,-13738.,-1689.8,-1331.9,-5205.5,-2799.2,-5723.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1410.000000000,6718.8,1729.3,1844.5,1609.8,2036.1,1406.5,2795.6,456.78,1932.4,390.12,700.93,762.27,0.0000,-3648.6,-6658.8,-304.34,-2717.2,-2549.4,-13738.,-1706.6,-1348.5,-5218.3,-2800.6,-5733.7,0.13340E+06,59628.,45676.,42869.,83103.,28637.,0.10265E+06,29663.,45347.,13536.,19453.,23432.,0.0000,-136.60,-141.36,-21.596,-129.49,-84.586,-524.53,-423.46,-43.193,-379.85,-45.993,-515.73
1411.000000000,6704.3,1720.0,1855.1,1602.3,2038.3,1404.2,2779.3,454.77,1939.5,389.54,699.95,762.90,0.0000,-3665.0,-6675.0,-306.76,-2716.2,-2557.9,-13739.,-1702.0,-1359.1,-5222.0,-2800.9,-5737.3,4105.2,1834.9,1405.6,1319.2,2557.4,881.25,3158.8,912.82,1395.5,416.53,598.63,721.09,0.0000,-4.2117,-4.3531,-0.66459,-3.9886,-2.6053,-16.142,-13.031,-1.3292,-11.689,-1.4154,-15.870
1412.000000000,6597.5,1702.1,1851.3,1587.0,2033.8,1415.1,2780.2,457.25,1901.0,390.20,702.80,764.40,0.0000,-3633.6,-6667.1,-304.78,-2715.5,-2537.5,-13739.,-1697.7,-1344.6,-5210.8,-2798.6,-5729.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1413.000000000,6573.1,1712.9,1849.4,1572.7,2090.4,1424.2,2796.6,456.22,1904.9,389.25,710.96,763.24,0.0000,-3624.2,-6657.0,-302.64,-2714.7,-2533.5,-13741.,-1694.4,-1337.5,-5206.5,-2798.0,-5725.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1414.000000000,6462.7,1704.7,1828.7,1560.2,2105.6,1410.2,2782.7,455.42,1908.9,390.27,706.83,767.78,0.0000,-3616.8,-6647.7,-300.98,-2713.6,-2530.4,-13743.,-1692.0,-1332.8,-5204.2,-2797.5,-5723.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1415.000000000,6352.9,1668.9,1810.7,1569.5,2083.7,1390.1,2763.9,448.46,1920.1,393.48,709.69,782.15,0.0000,-3609.6,-6638.9,-299.71,-2712.3,-2527.2,-13743.,-1690.2,-1329.2,-5203.0,-2796.8,-5721.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1416.000000000,6411.2,1679.5,1796.6,1600.6,2096.3,1410.8,2768.6,443.79,1942.6,394.83,704.14,790.99,0.0000,-3602.9,-6630.1,-298.72,-2710.9,-2524.3,-13741.,-1689.0,-1326.1,-5201.2,-2795.9,-5719.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1417.000000000,6495.8,1696.8,1793.0,1631.6,2092.0,1411.8,2751.7,440.57,1961.1,395.47,713.17,791.25,0.0000,-3597.2,-6622.5,-297.93,-2709.8,-2521.7,-13740.,-1688.1,-1323.3,-5199.9,-2795.8,-5718.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1418.000000000,6490.8,1709.9,1770.6,1645.3,2084.0,1404.7,2722.4,441.65,1964.7,393.28,710.11,796.53,0.0000,-3591.7,-6615.8,-297.28,-2708.5,-2519.1,-13739.,-1687.5,-1320.7,-5198.8,-2795.2,-5717.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1419.000000000,6490.0,1718.9,1760.2,1641.9,2084.4,1380.9,2703.3,438.44,1966.7,394.52,704.42,806.40,0.0000,-3586.2,-6609.3,-296.72,-2707.1,-2516.3,-13737.,-1687.0,-1318.3,-5197.8,-2794.5,-5716.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1420.000000000,6490.5,1710.9,1771.0,1644.6,2090.1,1374.7,2656.1,438.50,1964.6,391.32,698.33,813.05,0.0000,-3580.7,-6602.8,-296.23,-2705.7,-2513.6,-13736.,-1686.7,-1316.1,-5197.0,-2793.8,-5715.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1421.000000000,6583.1,1698.5,1787.1,1621.6,2119.8,1354.8,2641.2,434.77,1938.7,391.58,690.01,814.88,0.0000,-3575.4,-6596.3,-295.79,-2704.4,-2511.2,-13734.,-1686.4,-1314.1,-5196.2,-2793.2,-5715.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1422.000000000,6566.9,1713.3,1773.9,1636.8,2155.5,1351.0,2623.2,426.69,1924.8,396.30,701.17,811.12,0.0000,-3570.6,-6590.7,-295.39,-2703.2,-2508.8,-13732.,-1686.2,-1312.2,-5195.5,-2792.7,-5714.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1423.000000000,6544.8,1710.6,1768.3,1635.1,2189.1,1339.9,2660.9,426.76,1937.0,397.12,709.06,810.13,0.0000,-3565.9,-6586.2,-294.98,-2701.8,-2506.5,-13730.,-1686.0,-1310.6,-5195.1,-2792.4,-5714.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1424.000000000,6679.9,1710.3,1759.9,1641.5,2243.0,1329.2,2689.9,431.22,1969.2,392.21,716.02,810.16,0.0000,-3561.4,-6582.2,-294.61,-2700.4,-2504.2,-13729.,-1685.9,-1309.1,-5194.7,-2792.2,-5713.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1425.000000000,6878.6,1727.7,1776.2,1652.1,2263.3,1345.3,2738.3,434.50,1946.5,390.41,709.12,806.10,0.0000,-3557.0,-6578.6,-294.25,-2698.6,-2502.1,-13727.,-1685.7,-1307.7,-5194.3,-2791.7,-5713.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1426.000000000,7127.7,1756.2,1814.9,1646.9,2253.7,1378.8,2722.3,429.97,1956.4,394.62,708.78,804.84,0.0000,-3596.7,-6598.4,-297.90,-2697.0,-2527.9,-13727.,-1687.3,-1325.5,-5205.8,-2794.1,-5721.2,12074.,5396.9,4134.2,3880.1,7521.7,2591.9,9290.7,2684.8,4104.4,1225.1,1760.7,2120.8,0.0000,-12.267,-12.744,-1.9547,-11.666,-7.5740,-47.489,-38.304,-3.9094,-34.370,-4.1614,-46.639
1427.000000000,7375.5,1739.1,1837.5,1615.3,2275.6,1372.8,2706.7,430.79,1953.2,394.68,711.67,804.52,0.0000,-3571.3,-6597.5,-297.37,-2695.4,-2509.2,-13726.,-1686.8,-1317.8,-5197.8,-2792.6,-5715.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1428.000000000,7376.1,1762.0,1831.4,1627.9,2266.8,1377.5,2709.7,432.08,1964.0,397.63,717.24,802.88,0.0000,-3563.7,-6592.9,-296.31,-2693.9,-2504.9,-13724.,-1686.3,-1314.0,-5195.3,-2791.8,-5713.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1429.000000000,7360.0,1768.0,1833.4,1612.3,2276.9,1388.8,2702.5,433.55,1972.5,398.84,715.31,814.87,0.0000,-3558.5,-6587.7,-295.34,-2692.5,-2502.2,-13723.,-1686.0,-1311.5,-5194.0,-2791.1,-5712.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1430.000000000,7266.3,1771.6,1857.9,1612.1,2243.3,1392.0,2717.3,431.34,1965.2,401.61,696.31,829.41,0.0000,-3553.8,-6582.9,-294.53,-2691.0,-2499.9,-13722.,-1685.7,-1309.4,-5193.2,-2790.2,-5712.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1431.000000000,7237.3,1789.4,1865.8,1602.2,2236.9,1389.2,2727.0,429.50,1951.4,403.52,684.63,836.35,0.0000,-3549.5,-6578.8,-293.86,-2689.7,-2497.7,-13721.,-1685.4,-1307.6,-5192.5,-2789.5,-5711.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1432.000000000,7247.7,1803.6,1876.5,1585.3,2255.1,1398.4,2763.1,430.83,1955.1,406.16,684.58,833.83,0.0000,-3545.4,-6574.5,-293.28,-2688.3,-2495.6,-13720.,-1685.2,-1305.9,-5191.9,-2788.6,-5710.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1433.000000000,7483.5,1795.9,1893.5,1584.2,2260.6,1398.9,2751.5,429.85,1967.0,402.55,676.88,833.61,0.0000,-3585.2,-6593.3,-296.75,-2687.1,-2521.5,-13720.,-1691.9,-1323.2,-5204.2,-2790.2,-5719.2,50994.,22793.,17460.,16387.,31767.,10947.,39238.,11339.,17334.,5174.1,7436.1,8957.1,0.0000,-51.675,-53.742,-8.2554,-49.173,-31.808,-200.49,-161.68,-16.511,-145.11,-17.569,-196.79
1434.000000000,7584.4,1760.4,1820.6,1587.6,2259.4,1410.0,2745.4,424.44,1936.4,398.35,676.33,836.89,0.0000,-3603.8,-6614.6,-300.12,-2686.0,-2530.7,-13720.,-1701.7,-1335.2,-5210.4,-2790.6,-5725.3,86402.,38620.,29584.,27766.,53825.,18548.,66484.,19212.,29371.,8766.8,12599.,15177.,0.0000,-87.724,-91.111,-13.988,-83.364,-53.950,-339.67,-273.96,-27.975,-245.87,-29.769,-333.41
1435.000000000,7618.1,1773.6,1789.8,1585.2,2253.5,1407.1,2754.6,425.07,1922.1,399.38,678.23,837.87,0.0000,-3618.9,-6634.3,-302.81,-2685.0,-2537.5,-13721.,-1736.4,-1344.8,-5220.9,-2790.7,-5738.0,0.29054E+06,0.12986E+06,99480.,93365.,0.18099E+06,62369.,0.22356E+06,64603.,98763.,29479.,42367.,51033.,0.0000,-295.63,-306.62,-47.035,-280.50,-181.55,-1142.3,-921.55,-94.071,-826.77,-100.11,-1121.1
1436.000000000,7731.7,1896.0,1841.7,1565.9,2291.9,1527.5,2942.4,443.17,1937.9,424.93,720.13,891.42,0.0000,-3638.8,-6655.6,-305.03,-2686.4,-2550.7,-13727.,-1726.9,-1353.1,-5227.1,-2793.7,-5744.2,28524.,12750.,9766.7,9166.4,17769.,6123.2,21949.,6342.6,9696.3,2894.2,4159.5,5010.3,0.0000,-29.202,-30.169,-4.6178,-27.633,-17.992,-112.40,-90.560,-9.2356,-81.219,-9.8400,-110.24
1437.000000000,7732.3,1873.8,1851.7,1562.0,2289.9,1466.0,2875.4,429.05,1922.5,436.88,728.69,903.16,0.0000,-3611.9,-6653.0,-302.84,-2687.1,-2530.2,-13731.,-1715.3,-1338.2,-5220.3,-2794.5,-5736.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1438.000000000,7735.9,1860.0,1799.8,1583.9,2317.3,1396.2,2821.1,418.28,1912.0,429.42,729.84,897.48,0.0000,-3602.9,-6641.7,-300.54,-2687.5,-2523.8,-13732.,-1706.6,-1330.9,-5215.4,-2795.5,-5731.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1439.000000000,7752.5,1818.4,1812.3,1592.1,2349.9,1369.4,2823.8,428.24,1905.6,419.66,742.49,896.15,0.0000,-3595.3,-6631.8,-298.80,-2686.8,-2519.4,-13732.,-1700.2,-1326.2,-5211.7,-2797.2,-5727.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1440.000000000,7781.2,1813.5,1810.4,1598.5,2357.7,1386.1,2827.3,434.43,1949.5,417.54,753.34,893.14,0.0000,-3588.6,-6623.0,-297.54,-2685.5,-2516.5,-13733.,-1695.7,-1322.6,-5208.3,-2798.9,-5724.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1441.000000000,7806.7,1810.9,1799.6,1600.0,2354.4,1400.5,2834.4,439.31,1970.0,422.15,758.61,900.79,0.0000,-3582.8,-6616.3,-296.60,-2684.1,-2513.7,-13733.,-1692.6,-1319.6,-5205.7,-2800.9,-5721.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1442.000000000,7862.1,1795.4,1770.0,1606.5,2372.0,1403.0,2854.3,429.05,1976.4,425.47,747.04,906.47,0.0000,-3578.1,-6608.4,-295.85,-2682.7,-2510.7,-13733.,-1690.4,-1317.0,-5203.2,-2801.1,-5719.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1443.000000000,7817.5,1777.1,1756.3,1620.3,2398.9,1405.3,2880.1,447.13,1987.5,427.21,741.64,898.09,0.0000,-3618.0,-6623.6,-299.23,-2681.6,-2535.9,-13734.,-1689.9,-1334.8,-5212.7,-2802.3,-5726.2,6930.1,3097.6,2372.8,2227.0,4317.1,1487.7,5332.5,1540.9,2355.7,703.16,1010.6,1217.3,0.0000,-7.0690,-7.3207,-1.1219,-6.6974,-4.3438,-27.301,-22.013,-2.2438,-19.739,-2.3905,-26.804
1444.000000000,7764.6,1751.7,1751.1,1610.7,2416.5,1386.3,2827.8,440.22,1978.7,429.68,736.96,888.75,0.0000,-3591.9,-6619.0,-298.52,-2680.5,-2516.3,-13734.,-1688.6,-1325.4,-5203.8,-2800.0,-5720.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1445.000000000,7806.1,1741.2,1788.5,1596.3,2400.3,1385.6,2848.1,432.76,2002.1,422.62,733.91,883.05,0.0000,-3583.8,-6611.8,-297.34,-2679.4,-2511.5,-13734.,-1687.6,-1320.7,-5200.7,-2798.5,-5717.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1446.000000000,7921.7,1732.2,1772.9,1600.0,2403.5,1370.2,2812.1,432.80,1998.3,421.71,731.21,892.94,0.0000,-3578.1,-6604.6,-296.31,-2678.3,-2508.2,-13734.,-1687.1,-1317.7,-5199.1,-2797.4,-5716.5,1306.2,583.87,447.26,419.77,813.74,280.41,1005.1,290.45,444.03,132.54,190.48,229.44,0.0000,-1.3293,-1.3791,-0.21147,-1.2608,-0.81443,-5.1457,-4.1482,-0.42294,-3.7202,-0.45040,-5.0506
1447.000000000,7931.1,1734.9,1778.3,1574.6,2398.6,1369.7,2810.2,436.79,1969.4,426.19,726.39,883.90,0.0000,-3573.2,-6597.9,-295.47,-2677.4,-2505.4,-13733.,-1686.5,-1315.2,-5197.9,-2796.0,-5715.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1448.000000000,7953.5,1737.3,1786.4,1579.5,2387.5,1355.2,2843.6,432.07,1953.0,418.74,730.51,878.93,0.0000,-3568.7,-6591.7,-294.77,-2676.6,-2502.9,-13733.,-1686.0,-1313.0,-5197.1,-2794.6,-5715.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1449.000000000,8016.6,1761.2,1807.9,1610.6,2405.7,1342.4,2862.9,427.10,1944.7,414.96,737.01,878.15,0.0000,-3564.2,-6586.3,-294.17,-2675.8,-2500.5,-13733.,-1685.7,-1311.0,-5196.5,-2793.9,-5714.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1450.000000000,7977.1,1762.1,1760.3,1632.2,2359.8,1348.3,2885.8,433.56,1943.8,414.58,733.42,889.41,0.0000,-3560.0,-6581.6,-293.62,-2675.0,-2498.4,-13732.,-1685.4,-1309.2,-5196.4,-2793.2,-5714.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1451.000000000,8005.7,1758.9,1783.6,1616.2,2332.4,1369.2,2889.5,432.44,1956.3,416.88,732.29,893.35,0.0000,-3555.6,-6577.9,-293.11,-2674.5,-2496.2,-13731.,-1685.2,-1307.5,-5196.4,-2792.6,-5713.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1452.000000000,8063.5,1772.5,1789.1,1617.2,2343.5,1369.8,2904.2,431.41,1971.7,417.89,726.35,907.06,0.0000,-3595.3,-6597.9,-296.62,-2674.2,-2522.1,-13731.,-1686.0,-1325.3,-5207.8,-2794.6,-5721.5,6695.4,2992.7,2292.5,2151.6,4170.9,1437.3,5151.9,1488.8,2276.0,679.35,976.35,1176.1,0.0000,-6.7977,-7.0609,-1.0839,-6.4527,-4.1621,-26.374,-21.251,-2.1679,-19.064,-2.3075,-25.867
1453.000000000,8047.8,1783.5,1802.2,1604.1,2326.1,1353.0,2939.7,432.56,1952.9,421.43,725.02,905.89,0.0000,-3570.3,-6596.2,-295.99,-2674.0,-2503.4,-13730.,-1685.6,-1317.4,-5199.8,-2792.6,-5716.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1454.000000000,8070.8,1789.7,1845.7,1604.1,2595.7,1369.3,2965.7,429.74,1960.3,421.42,720.20,901.48,0.0000,-3607.3,-6614.9,-298.84,-2673.9,-2527.2,-13730.,-1687.0,-1333.5,-5209.7,-2794.0,-5722.5,11907.,5322.2,4076.9,3826.3,7417.5,2556.0,9162.0,2647.6,4047.5,1208.1,1736.3,2091.5,0.0000,-12.107,-12.562,-1.9276,-11.479,-7.4035,-46.903,-37.785,-3.8553,-33.899,-4.1033,-45.989
1455.000000000,8158.1,1770.4,1837.4,1598.4,2445.2,1355.6,2948.0,428.24,1955.3,421.95,716.71,891.81,0.0000,-3581.1,-6611.8,-297.62,-2674.0,-2507.9,-13729.,-1686.3,-1323.9,-5201.0,-2791.5,-5716.4,18.493,8.2662,6.3321,5.9429,11.521,3.9699,14.230,4.1122,6.2865,1.8764,2.6968,3.2484,0.0000,-0.18797E-01,-0.19512E-01,-0.29939E-02,-0.17826E-01,-0.11482E-01,-0.72848E-01,-0.58681E-01,-0.59878E-02,-0.52648E-01,-0.63727E-02,-0.71418E-01
1456.000000000,8204.7,1787.9,1837.3,1583.4,2421.7,1357.6,2933.9,422.92,1957.4,421.89,715.07,882.13,0.0000,-3573.2,-6605.5,-296.06,-2674.0,-2503.4,-13728.,-1685.8,-1318.9,-5198.3,-2790.1,-5714.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1457.000000000,8287.4,1801.2,1814.5,1578.7,2428.0,1349.9,2918.9,418.40,1985.3,416.94,716.40,885.97,0.0000,-3567.9,-6599.1,-294.75,-2674.2,-2500.7,-13727.,-1685.3,-1315.5,-5197.0,-2788.9,-5712.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1458.000000000,8507.8,1770.0,1830.5,1580.9,2389.4,1371.9,2908.4,417.24,2021.2,420.22,717.25,885.76,0.0000,-3563.3,-6593.2,-293.72,-2674.3,-2498.9,-13726.,-1685.0,-1312.8,-5196.1,-2788.3,-5711.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1459.000000000,8567.7,1755.7,1808.0,1611.1,2397.1,1368.9,2921.2,416.70,2013.4,418.01,719.37,892.77,0.0000,-3559.0,-6587.7,-292.91,-2674.0,-2497.2,-13725.,-1684.7,-1310.4,-5195.6,-2787.6,-5711.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1460.000000000,8605.8,1742.7,1807.2,1618.3,2399.7,1384.6,2946.1,415.08,2030.1,416.89,724.66,887.89,0.0000,-3598.7,-6605.6,-296.24,-2673.7,-2523.3,-13724.,-1685.0,-1327.6,-5206.5,-2789.7,-5718.6,2952.2,1319.6,1010.8,948.68,1839.1,633.73,2271.6,656.43,1003.5,299.54,430.49,518.55,0.0000,-2.9974,-3.1122,-0.47793,-2.8434,-1.8308,-11.629,-9.3629,-0.95585,-8.4023,-1.0171,-11.393
1461.000000000,8586.9,1748.4,1801.4,1629.0,2406.0,1366.2,2950.0,412.37,2000.6,415.57,731.97,891.13,0.0000,-3573.1,-6602.5,-295.52,-2673.1,-2504.7,-13722.,-1684.8,-1318.9,-5198.3,-2787.8,-5712.9,468.84,209.56,160.53,150.66,292.07,100.64,360.76,104.25,159.37,47.571,68.368,82.353,0.0000,-0.47581,-0.49424,-0.75901E-01,-0.45150,-0.29040,-1.8467,-1.4868,-0.15180,-1.3343,-0.16152,-1.8092
1462.000000000,8468.9,1736.1,1799.2,1632.2,2409.3,1379.3,3014.0,411.87,1972.1,416.67,733.70,887.12,0.0000,-3565.1,-6596.2,-294.33,-2672.5,-2500.6,-13721.,-1684.5,-1314.3,-5195.8,-2786.8,-5711.1,74.548,33.321,25.525,23.956,46.440,16.003,57.362,16.576,25.341,7.5640,10.871,13.094,0.0000,-0.75606E-01,-0.78569E-01,-0.12069E-01,-0.71771E-01,-0.46134E-01,-0.29365,-0.23639,-0.24137E-01,-0.21215,-0.25682E-01,-0.28763
1463.000000000,8577.8,1725.5,1799.5,1649.4,2430.0,1382.4,3037.9,417.67,1967.1,416.35,740.26,889.20,0.0000,-3603.4,-6613.1,-297.29,-2672.0,-2525.9,-13721.,-1685.3,-1330.9,-5206.1,-2788.6,-5718.5,7147.2,3194.7,2447.2,2296.8,4452.4,1534.3,5499.6,1589.2,2429.6,725.19,1042.2,1255.4,0.0000,-7.2617,-7.5353,-1.1571,-6.8849,-4.4316,-28.155,-22.662,-2.3141,-20.339,-2.4624,-27.573
1464.000000000,8563.5,1727.7,1777.0,1644.3,2413.5,1368.3,3034.9,420.33,1928.1,413.36,736.92,890.20,0.0000,-3577.0,-6609.0,-296.27,-2671.3,-2506.8,-13720.,-1684.9,-1321.4,-5197.5,-2786.5,-5712.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1465.000000000,8536.0,1722.4,1778.0,1633.1,2404.5,1340.9,3007.8,419.08,1932.1,414.27,738.91,893.11,0.0000,-3568.3,-6601.6,-294.87,-2670.7,-2502.4,-13718.,-1684.6,-1316.5,-5194.8,-2785.3,-5710.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1466.000000000,8567.1,1707.7,1757.6,1624.2,2420.3,1319.0,2964.6,423.40,1937.5,415.37,739.38,897.26,0.0000,-3562.0,-6593.9,-293.69,-2670.1,-2499.5,-13717.,-1684.3,-1313.0,-5193.5,-2784.4,-5709.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1467.000000000,8590.5,1699.3,1749.4,1623.0,2427.6,1321.0,2960.3,425.16,1936.3,418.16,738.56,898.57,0.0000,-3556.5,-6586.9,-292.74,-2669.4,-2497.1,-13716.,-1684.1,-1310.3,-5192.6,-2783.6,-5709.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1468.000000000,8386.0,1684.2,1793.0,1622.1,2449.7,1314.0,2964.7,420.80,1921.3,415.73,741.35,898.88,0.0000,-3551.4,-6581.6,-291.97,-2668.6,-2494.8,-13715.,-1683.9,-1308.1,-5191.9,-2782.8,-5708.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1469.000000000,8358.5,1679.0,1793.9,1643.2,2465.8,1306.4,3011.4,422.39,1908.1,416.34,732.46,897.37,0.0000,-3546.7,-6577.3,-291.33,-2667.8,-2492.6,-13714.,-1683.7,-1306.1,-5191.3,-2781.9,-5707.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1470.000000000,8670.4,1662.4,1758.6,1660.1,2318.9,1316.7,3019.1,430.93,1900.5,412.57,738.99,886.90,0.0000,-3542.3,-6573.3,-290.77,-2667.1,-2490.6,-13714.,-1683.6,-1304.3,-5190.8,-2781.0,-5707.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1471.000000000,8728.2,1633.2,1749.1,1659.7,2327.3,1318.2,3022.5,432.58,1909.5,407.52,741.19,889.38,0.0000,-3538.1,-6569.5,-290.29,-2666.4,-2488.5,-13712.,-1683.4,-1302.7,-5190.4,-2780.1,-5706.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1472.000000000,8767.3,1625.1,1730.8,1660.1,2322.8,1302.8,2989.7,439.12,1917.9,409.15,744.45,889.41,0.0000,-3534.1,-6565.7,-289.84,-2665.8,-2486.5,-13711.,-1683.3,-1301.1,-5190.0,-2779.3,-5706.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1473.000000000,8729.4,1622.9,1734.0,1646.8,2477.2,1293.7,2973.9,437.71,1904.6,409.09,742.33,887.86,0.0000,-3530.2,-6562.1,-289.43,-2665.2,-2484.5,-13710.,-1683.2,-1299.6,-5189.6,-2778.5,-5705.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1474.000000000,8674.9,1611.2,1732.7,1658.5,2578.2,1281.4,2979.8,432.38,1915.5,405.78,740.81,884.77,0.0000,-3526.3,-6558.8,-289.06,-2664.5,-2482.5,-13709.,-1683.1,-1298.5,-5189.2,-2777.8,-5705.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1475.000000000,8678.0,1624.4,1743.0,1688.9,2568.4,1293.2,2999.8,426.70,1903.6,407.63,737.57,885.18,0.0000,-3566.0,-6578.9,-292.68,-2664.0,-2508.5,-13709.,-1684.6,-1315.4,-5200.5,-2779.8,-5713.5,11000.,4916.6,3766.2,3534.8,6852.3,2361.2,8463.8,2445.8,3739.1,1116.1,1604.0,1932.1,0.0000,-11.111,-11.562,-1.7807,-10.569,-6.7791,-43.343,-34.841,-3.5615,-31.286,-3.7881,-42.375
1476.000000000,8699.9,1645.4,1748.0,1712.0,2586.8,1286.3,3017.3,420.22,1891.2,407.82,734.96,889.51,0.0000,-3584.8,-6600.8,-296.17,-2663.4,-2517.8,-13708.,-1687.1,-1327.6,-5204.3,-2780.3,-5717.0,21768.,9729.8,7453.3,6995.2,13560.,4672.8,16750.,4840.2,7399.6,2208.7,3174.3,3823.6,0.0000,-22.024,-22.893,-3.5240,-20.931,-13.435,-85.774,-68.945,-7.0480,-61.912,-7.4970,-83.851
1477.000000000,8692.3,1646.1,1761.0,1706.0,2416.5,1279.0,3040.3,420.05,1905.3,409.20,733.84,888.92,0.0000,-3600.0,-6621.0,-298.96,-2662.9,-2524.8,-13707.,-1692.5,-1337.3,-5206.9,-2780.5,-5720.2,47893.,21407.,16398.,15391.,29835.,10281.,36852.,10649.,16280.,4859.5,6983.9,8412.5,0.0000,-48.545,-50.405,-7.7534,-46.087,-29.590,-188.71,-151.69,-15.507,-136.21,-16.495,-184.47
1478.000000000,8703.0,1633.2,1756.3,1693.4,2464.6,1260.6,3047.8,417.44,1893.3,408.74,731.12,897.43,0.0000,-3569.6,-6615.8,-297.15,-2662.2,-2503.1,-13705.,-1690.0,-1324.5,-5196.5,-2778.0,-5713.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1479.000000000,8700.3,1619.3,1768.3,1689.5,2471.6,1263.2,3067.0,416.43,1904.3,409.86,738.64,894.92,0.0000,-3603.5,-6630.0,-299.10,-2661.5,-2525.5,-13704.,-1696.2,-1338.6,-5206.0,-2779.3,-5721.1,61155.,27335.,20939.,19652.,38097.,13128.,47056.,13598.,20788.,6205.1,8917.7,10742.,0.0000,-62.071,-64.407,-9.9004,-58.879,-37.773,-240.97,-193.68,-19.801,-173.92,-21.061,-235.51
1480.000000000,8692.0,1614.6,1752.3,1688.8,2490.6,1246.7,3047.7,415.68,1878.9,408.69,747.18,900.33,0.0000,-3574.7,-6622.9,-297.26,-2660.9,-2505.3,-13702.,-1692.6,-1326.8,-5197.0,-2777.0,-5715.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1481.000000000,8568.9,1619.3,1744.7,1704.9,2497.0,1249.4,3032.3,412.71,1872.6,405.78,747.53,895.66,0.0000,-3564.4,-6612.9,-295.29,-2660.2,-2500.2,-13701.,-1689.7,-1320.7,-5193.4,-2775.8,-5713.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1482.000000000,8773.5,1617.6,1754.8,1711.8,2521.5,1263.1,3046.7,415.01,1862.4,403.66,749.86,896.82,0.0000,-3557.0,-6603.6,-293.72,-2659.6,-2497.1,-13700.,-1687.6,-1316.3,-5191.2,-2774.9,-5711.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1483.000000000,8773.2,1638.2,1748.4,1716.1,2541.8,1277.7,3074.0,413.95,1847.7,402.91,750.40,890.69,0.0000,-3550.9,-6595.4,-292.53,-2659.0,-2495.2,-13700.,-1686.1,-1312.9,-5189.7,-2774.5,-5710.1,0.27207,0.12161,0.93157E-01,0.87431E-01,0.16949,0.58405E-01,0.20935,0.60497E-01,0.92485E-01,0.27606E-01,0.39674E-01,0.47790E-01,0.0000,-0.27554E-03,-0.28640E-03,-0.44046E-04,-0.26177E-03,-0.16760E-03,-0.10725E-02,-0.86157E-03,-0.88092E-04,-0.77372E-03,-0.93686E-04,-0.10477E-02
1484.000000000,8746.2,1628.8,1738.9,1719.2,2540.2,1250.9,3060.3,418.89,1843.5,399.88,751.02,884.67,0.0000,-3545.9,-6588.7,-291.62,-2658.2,-2492.8,-13701.,-1685.0,-1310.0,-5188.5,-2773.9,-5709.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1485.000000000,8647.6,1621.4,1766.3,1717.9,2537.4,1234.4,3042.8,423.08,1847.7,401.94,751.41,878.18,0.0000,-3540.9,-6582.9,-290.89,-2657.3,-2490.4,-13700.,-1684.2,-1307.6,-5187.6,-2773.2,-5708.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1486.000000000,8677.8,1616.3,1798.5,1724.1,2523.8,1240.9,3037.5,428.89,1865.6,402.19,753.16,873.05,0.0000,-3536.1,-6577.6,-290.29,-2656.5,-2488.1,-13700.,-1683.7,-1305.7,-5187.2,-2772.7,-5707.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1487.000000000,8596.8,1623.7,1798.7,1728.0,2519.9,1249.6,3029.1,423.99,1877.1,399.56,758.04,873.72,0.0000,-3531.5,-6572.8,-289.77,-2655.7,-2485.7,-13699.,-1683.3,-1304.0,-5186.6,-2772.2,-5706.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1488.000000000,8533.8,1618.5,1792.0,1736.4,2495.1,1241.4,3006.6,419.38,1852.3,396.78,758.87,869.49,0.0000,-3526.9,-6568.2,-289.31,-2654.8,-2483.2,-13697.,-1682.9,-1302.3,-5186.0,-2771.5,-5705.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1489.000000000,8547.8,1618.5,1776.8,1723.5,2474.5,1239.6,3019.3,418.52,1833.1,396.22,763.05,870.03,0.0000,-3566.0,-6586.4,-292.88,-2654.3,-2508.7,-13696.,-1683.2,-1319.1,-5197.2,-2773.7,-5713.2,3484.0,1557.3,1192.9,1119.6,2170.3,747.89,2680.8,774.68,1184.3,353.50,508.04,611.96,0.0000,-3.5205,-3.6608,-0.56402,-3.3480,-2.1443,-13.731,-11.030,-1.1280,-9.9072,-1.1994,-13.412
1490.000000000,8645.6,1627.1,1770.1,1702.7,2467.1,1215.5,3022.2,419.58,1849.2,396.24,760.25,864.21,0.0000,-3540.3,-6583.6,-292.32,-2653.9,-2489.7,-13694.,-1682.9,-1311.2,-5188.9,-2771.9,-5707.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1491.000000000,8527.9,1652.0,1781.7,1693.2,2430.9,1201.1,3020.9,421.44,1882.2,394.12,751.54,862.67,0.0000,-3532.4,-6577.6,-291.25,-2653.4,-2485.3,-13691.,-1682.7,-1307.1,-5186.2,-2770.9,-5705.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1492.000000000,8635.5,1627.4,1779.9,1702.5,2408.9,1195.1,3013.1,423.24,1868.6,391.95,750.23,859.54,0.0000,-3526.7,-6571.6,-290.31,-2652.8,-2482.4,-13689.,-1682.4,-1304.4,-5185.0,-2770.2,-5705.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1493.000000000,8648.0,1612.8,1771.0,1690.3,2417.3,1201.5,2996.8,428.29,1841.3,387.93,747.71,856.07,0.0000,-3521.6,-6566.1,-289.54,-2652.0,-2480.0,-13687.,-1682.3,-1302.2,-5184.1,-2769.5,-5704.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1494.000000000,8611.6,1599.3,1788.6,1708.5,2422.8,1219.2,3002.2,425.85,1844.4,389.41,748.61,848.50,0.0000,-3517.0,-6561.5,-288.94,-2651.2,-2477.8,-13686.,-1682.1,-1300.3,-5183.5,-2769.0,-5704.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1495.000000000,8596.6,1610.1,1785.5,1723.9,2404.5,1213.8,3009.7,421.25,1870.1,389.60,751.48,848.26,0.0000,-3512.6,-6557.5,-288.44,-2650.4,-2475.6,-13684.,-1682.0,-1298.5,-5182.9,-2768.7,-5703.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1496.000000000,8467.6,1626.4,1785.2,1721.2,2384.9,1197.0,2995.7,421.68,1881.5,390.24,759.49,849.45,0.0000,-3508.4,-6553.3,-288.02,-2649.6,-2473.4,-13682.,-1681.9,-1297.0,-5182.4,-2768.3,-5703.4,29.222,13.062,10.006,9.3907,18.204,6.2731,22.486,6.4978,9.9336,2.9651,4.2613,5.1330,0.0000,-0.29403E-01,-0.30633E-01,-0.47308E-02,-0.28026E-01,-0.17867E-01,-0.11507,-0.92471E-01,-0.94617E-02,-0.83081E-01,-0.10056E-01,-0.11242
1497.000000000,8506.1,1620.5,1861.3,1752.7,2387.0,1224.7,2998.7,417.06,1885.4,390.20,755.01,850.75,0.0000,-3547.8,-6572.6,-291.62,-2649.2,-2499.2,-13681.,-1682.1,-1313.5,-5193.4,-2770.4,-5711.0,1924.0,859.99,658.77,618.28,1198.6,413.02,1480.4,427.81,654.02,195.22,280.56,337.95,0.0000,-1.9384,-2.0172,-0.31148,-1.8463,-1.1786,-7.5755,-6.0878,-0.62295,-5.4699,-0.66213,-7.4011
1498.000000000,8525.6,1600.8,1893.3,1755.3,2375.8,1194.5,3013.6,417.65,1873.5,388.30,749.50,841.95,0.0000,-3522.6,-6571.1,-291.10,-2648.8,-2480.6,-13679.,-1681.9,-1306.1,-5185.0,-2768.5,-5705.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1499.000000000,8553.3,1619.9,1907.9,1759.3,2367.4,1175.6,3030.1,415.27,1876.8,383.46,746.29,834.63,0.0000,-3515.2,-6566.4,-290.07,-2648.3,-2476.4,-13678.,-1681.8,-1302.4,-5182.3,-2767.7,-5703.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1500.000000000,8680.8,1608.5,1876.5,1760.3,2368.4,1169.4,3027.2,415.53,1880.1,377.74,744.39,828.67,0.0000,-3510.0,-6561.3,-289.15,-2647.8,-2473.6,-13676.,-1681.6,-1299.8,-5181.1,-2766.8,-5703.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1501.000000000,8569.0,1575.6,1850.6,1771.3,2385.9,1154.3,3025.5,414.70,1877.3,375.54,740.32,825.31,0.0000,-3505.5,-6555.9,-288.42,-2647.3,-2471.1,-13675.,-1681.5,-1297.7,-5180.4,-2765.8,-5702.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1502.000000000,8483.1,1574.5,1859.4,1785.1,2381.1,1150.3,3003.2,410.46,1879.7,376.12,736.30,819.94,0.0000,-3501.3,-6551.1,-287.82,-2646.6,-2468.8,-13673.,-1681.4,-1295.8,-5179.7,-2764.8,-5701.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1503.000000000,8436.1,1546.4,1867.5,1786.4,2371.4,1150.3,2978.8,408.84,1890.2,375.30,734.23,823.75,0.0000,-3497.0,-6546.7,-287.32,-2646.0,-2466.6,-13672.,-1681.3,-1294.2,-5178.9,-2763.9,-5701.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1504.000000000,8409.5,1550.1,1845.5,1801.9,2419.5,1148.2,2994.1,409.75,1909.2,371.68,735.58,825.22,0.0000,-3493.2,-6542.8,-286.89,-2645.4,-2464.4,-13670.,-1681.1,-1292.6,-5178.3,-2763.1,-5701.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1505.000000000,8217.3,1561.6,1845.7,1824.6,2440.3,1144.1,2989.4,409.28,1893.8,374.55,734.44,815.67,0.0000,-3489.3,-6539.3,-286.50,-2644.9,-2462.4,-13669.,-1681.1,-1291.2,-5177.7,-2762.4,-5700.7,67.282,30.074,23.037,21.621,41.913,14.443,51.771,14.961,22.871,6.8267,9.8112,11.818,0.0000,-0.67461E-01,-0.70344E-01,-0.10892E-01,-0.64416E-01,-0.40894E-01,-0.26467,-0.21276,-0.21785E-01,-0.19123,-0.23138E-01,-0.25857
1506.000000000,8324.2,1569.7,1842.2,1836.0,2425.6,1156.0,3004.4,411.14,1897.3,371.47,737.46,812.88,0.0000,-3528.6,-6559.2,-290.13,-2644.5,-2488.2,-13668.,-1707.4,-1307.2,-5194.1,-2764.2,-5715.3,0.19744E+06,88251.,67603.,63448.,0.12300E+06,42384.,0.15192E+06,43902.,67116.,20033.,28791.,34680.,0.0000,-198.23,-206.47,-31.964,-189.14,-120.23,-776.58,-624.44,-63.927,-561.15,-67.900,-758.73
1507.000000000,8375.9,1564.8,1828.6,1866.0,2437.7,1157.4,3019.9,410.34,1893.9,372.95,737.17,808.56,0.0000,-3503.7,-6557.8,-289.64,-2644.1,-2469.5,-13667.,-1700.7,-1300.2,-5188.6,-2762.2,-5713.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1508.000000000,8328.3,1564.2,1843.5,1859.8,2505.8,1173.0,3045.1,408.01,1896.4,375.04,737.05,814.23,0.0000,-3496.3,-6553.3,-288.63,-2643.8,-2465.7,-13666.,-1695.2,-1296.6,-5186.0,-2761.1,-5711.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1509.000000000,8316.9,1577.8,1854.5,1875.1,2494.1,1224.7,3059.4,413.36,1895.7,374.95,741.65,814.25,0.0000,-3535.5,-6571.9,-291.75,-2644.1,-2492.6,-13666.,-1691.5,-1312.3,-5195.5,-2763.5,-5717.4,3643.9,1628.7,1247.7,1171.0,2270.0,782.22,2803.8,810.24,1238.7,369.72,531.36,640.05,0.0000,-3.6638,-3.8121,-0.58991,-3.4943,-2.2234,-14.339,-11.527,-1.1798,-10.358,-1.2533,-14.007
1510.000000000,8212.6,1572.8,1842.0,1859.6,2503.8,1214.2,3031.0,409.97,1899.5,369.48,750.67,809.24,0.0000,-3511.3,-6571.3,-290.89,-2644.1,-2474.0,-13666.,-1688.4,-1304.2,-5185.8,-2761.6,-5710.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1511.000000000,8209.5,1547.0,1830.1,1852.7,2486.3,1196.7,3003.5,408.81,1889.9,368.60,749.69,807.63,0.0000,-3503.6,-6565.5,-289.63,-2643.8,-2469.5,-13664.,-1686.1,-1300.0,-5182.3,-2760.7,-5706.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1512.000000000,8083.9,1552.7,1830.8,1858.8,2486.8,1210.4,3023.7,409.90,1902.5,368.46,749.50,809.25,0.0000,-3541.6,-6582.6,-292.54,-2643.7,-2494.6,-13663.,-1688.0,-1315.7,-5192.2,-2762.4,-5713.4,26082.,11658.,8930.6,8381.7,16248.,5599.0,20070.,5799.6,8866.2,2646.5,3803.4,4581.4,0.0000,-26.242,-27.288,-4.2225,-25.020,-15.919,-102.62,-82.516,-8.4450,-74.144,-8.9696,-100.27
1513.000000000,8021.4,1573.0,1819.9,1863.7,2509.6,1204.3,3005.1,409.58,1887.4,368.25,753.52,807.65,0.0000,-3515.9,-6578.6,-291.51,-2643.8,-2475.4,-13661.,-1686.1,-1306.9,-5183.3,-2760.5,-5707.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1514.000000000,7894.8,1576.7,1823.9,1875.8,2513.8,1192.3,2979.3,413.15,1872.1,361.97,750.53,809.11,0.0000,-3508.0,-6571.5,-290.13,-2644.1,-2471.0,-13660.,-1684.5,-1302.2,-5180.1,-2759.5,-5704.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1515.000000000,7893.3,1577.7,1827.1,1872.4,2515.4,1182.3,2949.5,413.27,1862.5,359.78,750.51,808.73,0.0000,-3502.5,-6564.5,-288.98,-2644.4,-2468.3,-13658.,-1683.4,-1299.0,-5178.4,-2758.7,-5702.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1516.000000000,7901.4,1574.8,1834.3,1888.0,2506.6,1173.5,2936.1,411.26,1867.9,357.73,750.06,807.92,0.0000,-3497.8,-6558.2,-288.08,-2644.4,-2465.7,-13657.,-1682.6,-1296.3,-5177.2,-2758.2,-5701.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1517.000000000,7885.3,1576.0,1834.0,1894.1,2510.3,1168.9,2927.7,406.84,1867.9,355.74,742.56,802.74,0.0000,-3493.1,-6553.0,-287.37,-2644.4,-2463.0,-13656.,-1681.9,-1294.1,-5176.2,-2757.6,-5700.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1518.000000000,7929.0,1588.0,1845.8,1884.7,2524.4,1171.8,2941.1,404.76,1879.6,358.87,746.34,811.28,0.0000,-3488.4,-6548.0,-286.80,-2644.3,-2460.6,-13654.,-1681.5,-1292.1,-5175.5,-2757.2,-5699.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1519.000000000,7890.6,1592.1,1849.0,1875.3,2529.5,1175.9,2955.1,404.89,1865.2,358.39,741.75,817.96,0.0000,-3484.1,-6543.0,-286.33,-2644.2,-2458.4,-13653.,-1681.1,-1290.3,-5174.7,-2756.9,-5698.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1520.000000000,7879.9,1611.1,1862.9,1882.6,2528.8,1173.5,2966.6,405.11,1846.2,358.49,744.19,816.69,0.0000,-3480.2,-6538.8,-285.93,-2644.1,-2456.3,-13652.,-1680.9,-1288.7,-5173.8,-2756.7,-5697.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1521.000000000,7859.6,1603.3,1861.5,1894.1,2513.0,1170.8,2949.7,405.34,1842.5,361.52,741.50,808.59,0.0000,-3476.5,-6535.3,-285.57,-2644.0,-2454.4,-13651.,-1680.7,-1287.2,-5172.9,-2756.7,-5696.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1522.000000000,7859.3,1620.9,1868.9,1898.2,2500.9,1169.6,2943.9,405.68,1831.1,360.18,740.86,808.41,0.0000,-3473.3,-6532.2,-285.25,-2643.9,-2452.5,-13649.,-1680.5,-1285.8,-5172.3,-2756.5,-5696.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1523.000000000,7876.6,1615.8,1926.1,1894.3,2607.5,1166.3,2920.8,405.88,1815.4,359.19,738.76,810.47,0.0000,-3470.1,-6529.2,-284.94,-2643.6,-2450.7,-13648.,-1680.3,-1284.5,-5171.6,-2756.0,-5695.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1524.000000000,7869.4,1634.8,1900.3,1902.6,2733.1,1161.1,2903.1,404.86,1812.7,358.71,735.36,810.42,0.0000,-3466.9,-6526.5,-284.64,-2643.1,-2448.9,-13647.,-1680.2,-1283.3,-5170.9,-2755.5,-5695.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1525.000000000,7876.7,1646.5,1903.4,1915.6,2725.1,1177.3,2918.2,404.98,1815.2,361.48,734.20,808.48,0.0000,-3507.1,-6547.1,-288.34,-2642.8,-2475.0,-13647.,-1682.0,-1298.9,-5182.1,-2757.6,-5702.9,13412.,5995.1,4592.4,4310.1,8355.3,2879.2,10320.,2982.3,4559.3,1360.9,1955.8,2355.9,0.0000,-13.416,-13.981,-2.1713,-12.831,-8.1116,-52.675,-42.400,-4.3427,-38.116,-4.6084,-51.504
1526.000000000,7873.4,1637.4,1903.0,1902.2,2718.3,1160.8,2922.4,403.13,1819.1,362.53,728.87,814.35,0.0000,-3483.3,-6546.6,-287.90,-2642.4,-2456.4,-13646.,-1681.4,-1292.4,-5173.8,-2755.8,-5697.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1527.000000000,8008.5,1636.2,1901.1,1893.5,2716.4,1138.5,2930.4,406.12,1798.9,366.00,721.30,814.09,0.0000,-3476.9,-6542.7,-286.93,-2641.9,-2452.2,-13645.,-1681.0,-1289.1,-5171.2,-2754.8,-5695.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1528.000000000,8040.3,1629.5,1901.5,1893.5,2712.9,1129.1,2933.9,407.68,1783.4,361.80,715.94,811.63,0.0000,-3472.6,-6538.3,-286.06,-2641.5,-2449.5,-13644.,-1680.6,-1286.8,-5170.0,-2753.8,-5694.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1529.000000000,8033.3,1635.7,2027.4,1885.6,2711.1,1129.2,2936.2,404.99,1779.7,358.78,715.92,803.88,0.0000,-3468.9,-6533.7,-285.34,-2641.1,-2447.2,-13643.,-1680.3,-1285.0,-5169.2,-2752.9,-5693.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1530.000000000,7932.3,1633.8,2041.2,1869.8,2687.2,1119.4,2929.9,402.58,1781.7,356.32,716.68,808.16,0.0000,-3465.7,-6529.8,-284.76,-2640.7,-2445.2,-13642.,-1680.0,-1283.4,-5168.5,-2751.9,-5693.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1531.000000000,7933.3,1631.2,2042.2,1871.4,2523.4,1141.6,2899.6,398.30,1808.9,355.86,710.32,814.95,0.0000,-3505.7,-6549.7,-288.23,-2640.4,-2470.9,-13643.,-1680.3,-1298.8,-5179.4,-2753.5,-5700.7,3374.5,1508.4,1155.4,1084.4,2102.2,724.40,2596.6,750.35,1147.1,342.40,492.09,592.74,0.0000,-3.3721,-3.5147,-0.54631,-3.2263,-2.0350,-13.242,-10.663,-1.0926,-9.5884,-1.1589,-12.950
1532.000000000,7983.4,1611.5,2055.7,1864.7,2541.0,1143.7,2914.7,391.50,1804.3,356.18,702.18,818.05,0.0000,-3481.5,-6548.8,-287.64,-2640.2,-2452.2,-13641.,-1680.1,-1291.8,-5171.0,-2751.0,-5695.2,131.95,58.981,45.181,42.404,82.201,28.326,101.53,29.341,44.855,13.389,19.242,23.178,0.0000,-0.13183,-0.13743,-0.21362E-01,-0.12614,-0.79471E-01,-0.51771,-0.41692,-0.42724E-01,-0.37492,-0.45311E-01,-0.50632
1533.000000000,8011.8,1604.7,2070.8,1849.3,2545.3,1141.2,2900.3,392.07,1810.6,355.46,698.77,815.55,0.0000,-3474.8,-6544.0,-286.55,-2640.0,-2448.0,-13641.,-1679.9,-1288.1,-5168.5,-2749.5,-5693.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1534.000000000,8024.2,1595.3,2098.9,1835.3,2554.5,1135.1,2911.9,390.42,1806.3,355.44,699.00,812.28,0.0000,-3470.4,-6538.9,-285.60,-2639.8,-2445.4,-13640.,-1679.7,-1285.6,-5167.3,-2748.3,-5692.3,231.80,103.61,79.369,74.490,144.40,49.760,178.36,51.543,78.796,23.520,33.802,40.716,0.0000,-0.23135,-0.24131,-0.37527E-01,-0.22147,-0.13937,-0.90917,-0.73228,-0.75053E-01,-0.65858,-0.79580E-01,-0.88925
1535.000000000,8059.2,1581.7,2086.9,1824.4,2539.5,1134.5,2912.4,389.17,1802.2,351.87,700.02,812.63,0.0000,-3466.3,-6534.1,-284.83,-2639.7,-2443.3,-13639.,-1679.5,-1283.6,-5166.6,-2747.7,-5691.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1536.000000000,8215.0,1589.0,2071.1,1810.7,2533.7,1134.4,2910.2,387.51,1786.5,351.28,695.04,814.91,0.0000,-3462.5,-6529.8,-284.22,-2639.6,-2441.4,-13638.,-1679.3,-1281.9,-5166.1,-2747.1,-5691.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1537.000000000,8282.2,1583.5,2067.0,1817.0,2528.0,1116.0,2909.5,388.06,1803.4,352.51,692.12,812.21,0.0000,-3458.9,-6526.2,-283.71,-2639.4,-2439.6,-13638.,-1679.2,-1280.4,-5165.7,-2746.5,-5690.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1538.000000000,8166.5,1569.3,2065.7,1800.6,2548.8,1108.4,2910.3,388.40,1818.5,352.99,687.17,811.79,0.0000,-3455.5,-6523.1,-283.28,-2639.2,-2437.8,-13637.,-1679.1,-1279.1,-5165.3,-2745.9,-5690.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1539.000000000,8140.6,1559.7,2068.0,1790.1,2555.4,1112.3,2908.2,385.26,1819.9,351.73,680.74,819.10,0.0000,-3452.1,-6520.2,-282.90,-2638.9,-2436.1,-13636.,-1679.0,-1278.1,-5164.9,-2745.3,-5690.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1540.000000000,8178.5,1560.4,2081.8,1786.3,2546.6,1112.2,2903.7,378.80,1821.6,350.86,671.49,823.26,0.0000,-3449.2,-6517.4,-282.56,-2638.7,-2434.4,-13635.,-1678.9,-1277.1,-5164.4,-2744.7,-5689.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1541.000000000,8198.0,1574.5,2083.1,1785.5,2545.9,1105.9,2902.4,377.94,1813.1,350.33,668.46,821.28,0.0000,-3446.4,-6514.7,-282.24,-2638.4,-2432.7,-13634.,-1678.8,-1276.1,-5164.1,-2744.2,-5689.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1542.000000000,7993.2,1561.2,2084.5,1790.1,2550.3,1096.4,2906.7,378.05,1815.1,350.33,670.38,824.01,0.0000,-3443.7,-6512.5,-281.96,-2638.2,-2431.1,-13633.,-1678.7,-1275.2,-5163.8,-2743.8,-5689.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1543.000000000,7989.9,1556.0,2082.8,1779.5,2553.6,1090.1,2877.4,376.23,1824.7,350.37,665.71,820.70,0.0000,-3440.9,-6510.5,-281.71,-2638.1,-2429.6,-13632.,-1678.6,-1274.3,-5163.5,-2743.2,-5688.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1544.000000000,8199.0,1561.6,2081.5,1770.5,2576.7,1106.0,2873.1,376.04,1844.6,353.09,663.57,816.95,0.0000,-3481.0,-6531.5,-285.43,-2638.2,-2455.4,-13632.,-1678.9,-1289.0,-5174.7,-2745.3,-5696.6,2353.1,1051.8,805.71,756.18,1465.9,505.14,1810.6,523.23,799.90,238.76,343.14,413.33,0.0000,-2.3408,-2.4435,-0.38095,-2.2446,-1.4115,-9.2171,-7.4282,-0.76190,-6.6835,-0.80730,-9.0181
1545.000000000,8215.2,1551.3,2059.6,1773.0,2578.5,1090.5,2865.7,378.63,1872.8,353.43,667.65,814.52,0.0000,-3457.0,-6530.9,-285.03,-2638.3,-2437.3,-13630.,-1678.8,-1283.3,-5166.5,-2743.4,-5691.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1546.000000000,8291.2,1540.5,2051.9,1765.9,2578.5,1093.1,2864.4,371.58,1871.3,353.20,669.87,813.64,0.0000,-3451.0,-6527.0,-284.10,-2638.3,-2433.7,-13629.,-1678.6,-1280.4,-5164.0,-2742.5,-5689.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1547.000000000,8178.3,1552.0,2051.4,1754.8,2564.7,1093.6,2859.0,368.32,1858.5,351.80,667.79,812.88,0.0000,-3447.1,-6522.7,-283.27,-2638.2,-2431.6,-13628.,-1678.5,-1278.3,-5162.9,-2741.8,-5688.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1548.000000000,8051.7,1577.3,2044.1,1749.5,2545.5,1086.9,2847.3,366.00,1861.1,350.41,671.09,813.74,0.0000,-3443.9,-6518.7,-282.61,-2638.1,-2429.8,-13627.,-1678.3,-1276.6,-5162.1,-2741.2,-5687.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1549.000000000,8184.2,1601.0,2049.8,1755.7,2558.8,1090.3,2880.5,363.04,1852.1,347.80,668.51,815.62,0.0000,-3483.7,-6538.2,-286.06,-2638.3,-2455.6,-13627.,-1689.9,-1291.2,-5175.4,-2743.2,-5698.1,87363.,39050.,29913.,28074.,54423.,18754.,67223.,19426.,29697.,8864.3,12740.,15345.,0.0000,-86.913,-90.676,-14.143,-83.332,-52.346,-342.00,-275.71,-28.287,-248.10,-29.963,-334.66
1550.000000000,8174.1,1613.8,2038.8,1751.3,2549.7,1082.9,2883.2,362.59,1830.3,346.90,662.38,811.17,0.0000,-3459.6,-6536.9,-285.47,-2638.4,-2437.5,-13625.,-1686.9,-1284.8,-5168.1,-2741.4,-5694.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1551.000000000,8206.4,1606.5,1929.2,1743.1,2543.0,1077.6,2874.3,359.90,1833.3,347.42,657.10,815.96,0.0000,-3453.3,-6532.0,-284.41,-2638.3,-2433.8,-13624.,-1684.4,-1281.4,-5165.5,-2740.3,-5692.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1552.000000000,8328.2,1596.6,1930.4,1739.4,2547.7,1086.4,2871.6,358.51,1839.2,345.33,650.67,824.27,0.0000,-3449.2,-6526.8,-283.50,-2638.2,-2431.6,-13624.,-1682.5,-1279.0,-5163.9,-2739.2,-5690.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1553.000000000,8320.3,1591.6,1936.1,1744.3,2561.1,1090.1,2854.0,367.53,1837.9,341.91,648.30,818.79,0.0000,-3488.6,-6544.9,-286.76,-2638.0,-2457.2,-13624.,-1703.4,-1293.7,-5178.5,-2740.9,-5703.1,0.16659E+06,74464.,57042.,53535.,0.10378E+06,35762.,0.12819E+06,37043.,56630.,16903.,24293.,29262.,0.0000,-165.83,-172.89,-26.970,-158.92,-99.721,-651.94,-525.78,-53.940,-473.07,-57.124,-637.99
1554.000000000,8354.7,1602.6,1926.6,1747.6,2564.9,1070.2,2881.8,371.63,1809.4,342.24,647.69,820.04,0.0000,-3464.3,-6542.1,-286.05,-2637.8,-2438.7,-13623.,-1696.8,-1286.8,-5171.4,-2738.7,-5699.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1555.000000000,8632.1,1622.1,1943.9,1734.5,2582.6,1103.4,2916.7,377.95,1786.8,346.59,659.32,829.87,0.0000,-3458.6,-6535.7,-284.94,-2638.2,-2437.1,-13623.,-1691.5,-1283.2,-5168.4,-2738.3,-5696.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1556.000000000,8666.9,1626.9,1926.8,1718.6,2580.5,1078.7,2912.7,373.24,1776.7,341.87,671.92,825.44,0.0000,-3456.2,-6531.5,-284.02,-2638.3,-2435.7,-13624.,-1687.5,-1280.4,-5166.5,-2738.2,-5694.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1557.000000000,8658.9,1608.2,1904.3,1718.4,2584.8,1071.6,2899.7,373.71,1766.8,341.23,669.49,823.13,0.0000,-3453.5,-6526.7,-283.32,-2638.1,-2434.0,-13625.,-1684.7,-1278.3,-5165.5,-2737.9,-5692.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1558.000000000,8685.2,1589.9,1889.1,1724.9,2574.4,1066.5,2861.9,371.13,1748.4,339.43,667.41,822.36,0.0000,-3449.7,-6521.6,-282.77,-2637.8,-2431.5,-13624.,-1682.6,-1276.5,-5164.3,-2737.7,-5690.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1559.000000000,8716.2,1611.2,1871.5,1711.1,2577.8,1074.5,2867.3,368.65,1748.2,334.64,667.15,826.02,0.0000,-3446.6,-6516.3,-282.32,-2637.8,-2429.3,-13623.,-1681.2,-1275.0,-5162.9,-2737.6,-5688.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1560.000000000,8716.1,1604.3,1861.1,1706.9,2587.6,1066.8,2863.5,366.46,1746.7,328.99,665.52,821.25,0.0000,-3443.4,-6511.7,-281.95,-2637.6,-2427.4,-13622.,-1680.2,-1273.7,-5161.4,-2737.0,-5687.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1561.000000000,8702.4,1594.5,1849.6,1700.6,2577.9,1053.2,2849.9,367.09,1739.9,322.06,664.89,813.08,0.0000,-3440.4,-6507.9,-281.65,-2637.0,-2425.6,-13622.,-1679.5,-1272.5,-5160.2,-2736.9,-5686.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1562.000000000,8716.6,1601.8,1884.6,1707.7,2572.3,1068.5,2855.1,371.33,1742.9,321.17,668.03,807.97,0.0000,-3480.3,-6528.6,-285.39,-2636.3,-2451.2,-13622.,-1686.2,-1287.2,-5172.4,-2739.2,-5695.5,54074.,24170.,18515.,17377.,33686.,11608.,41608.,12024.,18381.,5486.7,7885.3,9498.2,0.0000,-53.801,-56.043,-8.7541,-51.585,-32.382,-211.67,-170.76,-17.508,-153.61,-18.540,-207.27
1563.000000000,8584.0,1611.8,1880.4,1708.9,2545.2,1064.4,2854.9,376.38,1759.8,318.76,664.27,795.24,0.0000,-3499.6,-6550.1,-288.99,-2635.8,-2460.5,-13622.,-1686.1,-1298.6,-5176.4,-2740.1,-5699.1,14994.,6702.2,5134.1,4818.5,9340.9,3218.8,11538.,3334.1,5097.1,1521.4,2186.5,2633.8,0.0000,-14.946,-15.550,-2.4275,-14.316,-8.9926,-58.690,-47.352,-4.8549,-42.596,-5.1413,-57.473
1564.000000000,8547.8,1624.8,1859.4,1716.7,2552.3,1059.4,2857.4,374.58,1739.0,318.54,661.76,797.46,0.0000,-3515.3,-6570.2,-291.87,-2635.5,-2467.4,-13621.,-1686.3,-1308.1,-5177.9,-2740.6,-5700.7,17524.,7832.7,6000.0,5631.2,10916.,3761.7,13484.,3896.5,5956.8,1778.0,2555.3,3078.0,0.0000,-17.500,-18.187,-2.8369,-16.744,-10.520,-68.582,-55.339,-5.6738,-49.781,-6.0086,-67.165
1565.000000000,8411.4,1628.1,1852.3,1718.2,2558.7,1057.1,2835.3,372.55,1759.7,319.94,662.24,797.60,0.0000,-3529.4,-6588.6,-294.14,-2635.1,-2473.3,-13621.,-1693.9,-1316.4,-5180.0,-2740.9,-5703.6,74386.,33249.,25470.,23904.,46339.,15968.,57238.,16540.,25286.,7547.6,10847.,13066.,0.0000,-74.418,-77.264,-12.042,-71.127,-44.674,-291.07,-234.92,-24.085,-211.31,-25.505,-285.09
1566.000000000,8439.4,1622.9,1833.7,1722.8,2585.0,1034.1,2837.8,373.70,1768.4,319.29,657.03,798.59,0.0000,-3498.8,-6581.4,-291.99,-2634.8,-2450.9,-13619.,-1689.6,-1303.7,-5169.0,-2738.4,-5696.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1567.000000000,8460.7,1628.2,1856.3,1729.9,2583.4,1030.7,2841.6,375.59,1783.6,322.08,655.18,800.34,0.0000,-3532.4,-6593.5,-293.70,-2634.6,-2473.1,-13620.,-1686.9,-1316.8,-5176.4,-2739.8,-5701.5,5115.3,2286.4,1751.5,1643.8,3186.6,1098.1,3936.0,1137.4,1738.8,519.02,745.92,898.50,0.0000,-5.1244,-5.3182,-0.82811,-4.8939,-3.0684,-20.014,-16.154,-1.6562,-14.531,-1.7536,-19.604
1568.000000000,8467.7,1647.2,1866.8,1735.1,2588.0,1059.8,2858.6,378.55,1786.4,323.28,660.68,805.89,0.0000,-3548.4,-6608.0,-295.74,-2634.9,-2481.9,-13620.,-1687.7,-1325.8,-5178.2,-2740.5,-5703.1,25277.,11298.,8654.8,8122.8,15746.,5426.1,19450.,5620.5,8592.4,2564.7,3686.0,4439.9,0.0000,-25.377,-26.305,-4.0921,-24.212,-15.202,-98.924,-79.836,-8.1842,-71.811,-8.6665,-96.886
1569.000000000,8539.5,1638.5,1857.9,1730.7,2584.7,1055.8,2849.6,377.19,1769.6,321.06,668.71,807.69,0.0000,-3518.9,-6599.6,-293.55,-2634.8,-2460.6,-13619.,-1684.9,-1312.1,-5166.7,-2738.3,-5695.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1570.000000000,8482.9,1623.4,1844.8,1743.0,2579.1,1045.7,2816.2,374.70,1765.2,318.35,673.34,802.60,0.0000,-3508.9,-6588.0,-291.27,-2634.3,-2454.6,-13619.,-1682.8,-1305.0,-5163.0,-2737.3,-5691.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1571.000000000,8465.0,1626.0,1841.2,1739.5,2599.9,1063.1,2818.3,376.29,1751.1,315.98,670.38,806.55,0.0000,-3501.8,-6576.6,-289.49,-2633.7,-2450.7,-13619.,-1681.2,-1300.1,-5160.9,-2736.4,-5689.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1572.000000000,8449.5,1637.0,1842.4,1732.7,2610.3,1060.6,2820.5,371.51,1738.2,316.46,675.51,798.98,0.0000,-3495.7,-6566.5,-288.16,-2633.1,-2447.4,-13619.,-1680.1,-1296.3,-5159.4,-2735.5,-5687.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1573.000000000,8411.6,1632.1,1836.7,1733.0,2602.5,1062.6,2797.2,374.41,1733.4,316.82,674.84,795.65,0.0000,-3490.0,-6557.8,-287.14,-2632.5,-2444.1,-13619.,-1679.3,-1293.0,-5158.3,-2734.7,-5686.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1574.000000000,8400.6,1626.7,1827.8,1720.5,2613.5,1062.1,2818.7,376.58,1738.7,314.84,679.12,797.76,0.0000,-3484.8,-6549.6,-286.34,-2632.0,-2441.2,-13618.,-1678.7,-1290.2,-5157.5,-2734.0,-5685.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1575.000000000,8294.5,1626.2,1836.9,1693.7,2600.6,1060.9,2830.6,376.44,1760.8,315.22,676.01,799.11,0.0000,-3480.2,-6542.4,-285.70,-2631.6,-2438.8,-13618.,-1678.3,-1287.7,-5156.6,-2733.4,-5684.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1576.000000000,8098.6,1624.5,1828.9,1688.9,2598.7,1051.9,2816.3,377.00,1777.0,315.02,672.09,792.60,0.0000,-3476.2,-6536.5,-285.18,-2631.1,-2436.4,-13617.,-1677.9,-1285.5,-5155.8,-2733.1,-5683.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1577.000000000,8092.4,1628.7,1816.0,1669.4,2585.4,1054.3,2806.3,379.98,1782.9,313.29,669.64,796.68,0.0000,-3472.4,-6531.8,-284.74,-2630.5,-2434.0,-13616.,-1677.7,-1283.5,-5155.1,-2732.6,-5683.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1578.000000000,8085.0,1611.6,1807.1,1655.8,2544.2,1056.7,2799.2,379.08,1781.9,310.24,671.99,799.33,0.0000,-3468.3,-6527.1,-284.35,-2629.8,-2431.7,-13615.,-1677.5,-1281.7,-5154.7,-2732.2,-5682.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1579.000000000,8085.9,1604.1,1807.4,1662.6,2528.6,1054.5,2793.5,375.24,1787.2,312.26,674.00,799.85,0.0000,-3464.5,-6522.8,-284.00,-2629.1,-2429.5,-13614.,-1677.3,-1280.0,-5154.2,-2731.9,-5682.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1580.000000000,8025.7,1600.2,1826.3,1663.0,2540.1,1039.3,2802.6,375.59,1789.7,312.15,677.72,799.23,0.0000,-3460.9,-6519.0,-283.67,-2628.5,-2427.3,-13613.,-1677.2,-1278.5,-5153.7,-2731.5,-5681.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1581.000000000,8176.2,1593.4,1828.1,1655.0,2535.0,1024.1,2776.0,374.34,1772.8,311.26,676.03,796.85,0.0000,-3457.6,-6515.0,-283.35,-2628.0,-2425.3,-13612.,-1677.1,-1277.0,-5153.2,-2731.0,-5681.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1582.000000000,8173.6,1604.2,1849.7,1653.4,2537.1,1021.8,2794.9,372.24,1766.7,310.13,667.16,794.35,0.0000,-3454.4,-6511.3,-283.03,-2627.4,-2423.3,-13611.,-1676.9,-1275.6,-5152.6,-2730.2,-5681.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1583.000000000,8194.1,1599.9,1863.5,1660.3,2517.4,1029.0,2782.4,369.52,1751.1,310.82,668.05,791.81,0.0000,-3451.2,-6507.9,-282.72,-2626.7,-2421.2,-13610.,-1676.9,-1274.3,-5152.0,-2729.6,-5681.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1584.000000000,8196.4,1599.5,1874.2,1637.8,2508.8,1037.1,2796.8,367.34,1756.4,311.49,666.95,786.82,0.0000,-3448.1,-6504.5,-282.42,-2625.8,-2419.1,-13609.,-1676.8,-1273.1,-5151.6,-2729.0,-5680.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1585.000000000,8281.5,1603.6,1874.2,1638.7,2539.6,1053.2,2798.4,365.71,1733.8,313.36,665.69,786.45,0.0000,-3445.0,-6501.7,-282.13,-2624.9,-2417.2,-13609.,-1676.7,-1271.9,-5151.3,-2728.4,-5680.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1586.000000000,8292.8,1606.9,1882.8,1635.1,2517.5,1040.2,2787.4,368.80,1728.9,311.74,660.39,787.21,0.0000,-3441.7,-6498.8,-281.85,-2624.1,-2415.2,-13609.,-1676.6,-1270.7,-5151.2,-2727.8,-5680.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1587.000000000,8316.1,1598.1,1894.4,1645.8,2507.5,1030.5,2759.9,372.99,1726.3,309.36,663.01,781.21,0.0000,-3438.8,-6495.5,-281.56,-2623.3,-2413.4,-13608.,-1676.5,-1269.7,-5150.8,-2727.3,-5680.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1588.000000000,8492.7,1591.4,1876.2,1643.3,2507.2,1019.4,2731.8,374.96,1718.7,305.79,666.68,779.87,0.0000,-3435.6,-6492.6,-281.28,-2622.5,-2411.6,-13608.,-1676.4,-1268.8,-5150.4,-2726.9,-5680.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1589.000000000,8483.6,1604.9,1877.4,1646.3,2506.5,1026.3,2730.3,372.95,1708.0,303.38,665.62,784.08,0.0000,-3432.7,-6490.2,-281.00,-2621.8,-2409.8,-13607.,-1676.4,-1268.1,-5150.0,-2726.6,-5679.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1590.000000000,8511.5,1593.1,1850.9,1649.8,2399.5,1033.9,2738.7,374.25,1702.3,301.62,658.97,786.32,0.0000,-3430.0,-6487.9,-280.72,-2621.1,-2408.1,-13606.,-1676.3,-1267.5,-5149.4,-2726.1,-5679.6,69.480,31.056,23.790,22.328,43.283,14.915,53.463,15.449,23.618,7.0498,10.132,12.204,0.0000,-0.68871E-01,-0.71866E-01,-0.11248E-01,-0.66108E-01,-0.41127E-01,-0.27141,-0.21919,-0.22496E-01,-0.19733,-0.23773E-01,-0.26586
1591.000000000,8494.3,1580.8,1850.5,1656.2,2382.6,1032.3,2707.6,374.21,1671.9,298.29,660.09,780.93,0.0000,-3427.4,-6485.7,-280.44,-2620.4,-2406.5,-13606.,-1676.2,-1266.8,-5148.9,-2725.6,-5679.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1592.000000000,8529.4,1571.9,1865.9,1667.2,2380.7,1062.2,2721.5,374.56,1670.0,296.49,658.40,775.47,0.0000,-3467.3,-6506.6,-284.12,-2619.8,-2432.2,-13606.,-1685.4,-1280.8,-5161.8,-2727.7,-5689.4,68988.,30836.,23622.,22170.,42977.,14810.,53084.,15340.,23451.,6999.9,10060.,12118.,0.0000,-68.454,-71.364,-11.169,-65.662,-40.907,-269.45,-217.63,-22.337,-195.92,-23.603,-263.93
1593.000000000,8623.6,1577.4,1872.3,1659.8,2393.1,1070.0,2759.0,374.40,1653.1,294.88,658.20,772.86,0.0000,-3443.5,-6506.3,-283.69,-2619.4,-2414.0,-13605.,-1683.0,-1275.7,-5154.6,-2725.9,-5685.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1594.000000000,8622.4,1552.6,1793.0,1677.6,2396.0,1064.9,2795.6,380.65,1644.9,294.01,656.79,771.65,0.0000,-3437.1,-6502.5,-282.72,-2618.9,-2410.3,-13604.,-1681.1,-1273.1,-5152.3,-2725.0,-5683.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1595.000000000,8563.6,1544.4,1717.4,1689.9,2397.2,1055.6,2798.3,384.64,1630.6,297.99,657.93,769.57,0.0000,-3432.9,-6498.3,-281.81,-2618.5,-2408.1,-13603.,-1679.6,-1271.4,-5150.9,-2724.3,-5681.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1596.000000000,8536.6,1559.9,1699.9,1686.6,2398.0,1048.7,2846.8,384.56,1630.2,300.36,656.90,769.95,0.0000,-3429.5,-6494.5,-281.05,-2618.1,-2406.3,-13603.,-1678.4,-1270.1,-5149.8,-2723.7,-5680.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1597.000000000,8595.3,1559.7,1691.5,1681.4,2416.3,1055.8,2829.6,383.14,1622.2,301.11,661.12,777.89,0.0000,-3426.7,-6491.2,-280.41,-2617.6,-2404.7,-13602.,-1677.6,-1269.0,-5148.8,-2722.8,-5679.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1598.000000000,8604.1,1563.3,1711.4,1692.3,2428.5,1064.3,2827.9,382.95,1624.7,301.76,669.11,777.03,0.0000,-3466.8,-6512.0,-283.83,-2617.1,-2430.5,-13602.,-1677.3,-1282.9,-5159.3,-2724.4,-5687.0,1698.6,759.25,581.61,545.86,1058.2,364.64,1307.0,377.70,577.42,172.35,247.70,298.37,0.0000,-1.6849,-1.7563,-0.27499,-1.6159,-1.0053,-6.6318,-5.3564,-0.54999,-4.8232,-0.58092,-6.4949
1599.000000000,8643.0,1561.0,1691.9,1689.5,2397.6,1051.5,2821.4,384.28,1608.1,299.50,668.53,778.39,0.0000,-3443.2,-6511.3,-283.20,-2616.6,-2412.4,-13602.,-1676.9,-1277.4,-5150.6,-2722.3,-5681.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1600.000000000,8659.4,1580.3,1684.8,1663.9,2386.4,1057.9,2814.7,379.78,1589.1,295.34,668.27,771.64,0.0000,-3437.1,-6506.7,-282.08,-2616.1,-2408.7,-13601.,-1676.5,-1274.3,-5147.6,-2721.1,-5678.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1601.000000000,8699.7,1578.2,1666.3,1661.4,2412.8,1088.6,2833.2,379.77,1582.2,296.54,667.05,768.49,0.0000,-3475.9,-6525.0,-285.06,-2616.1,-2433.8,-13601.,-1694.3,-1288.0,-5161.4,-2722.6,-5690.3,0.13517E+06,60419.,46283.,43438.,84206.,29017.,0.10401E+06,30056.,45949.,13715.,19711.,23743.,0.0000,-134.23,-139.80,-21.883,-128.63,-79.999,-527.62,-426.23,-43.766,-383.79,-46.219,-516.72
1602.000000000,8677.0,1599.3,1728.6,1651.0,2415.0,1110.9,2834.6,387.46,1567.4,298.94,667.26,762.99,0.0000,-3494.1,-6545.3,-288.07,-2616.2,-2443.3,-13601.,-1690.8,-1298.5,-5166.0,-2723.1,-5694.8,8887.4,3972.5,3043.0,2856.0,5536.5,1907.8,6838.6,1976.2,3021.1,901.76,1296.0,1561.1,0.0000,-8.8418,-9.1978,-1.4388,-8.4639,-5.2685,-34.689,-28.025,-2.8776,-25.234,-3.0389,-33.973
1603.000000000,8615.4,1597.7,1803.6,1643.1,2387.3,1120.3,2832.2,385.57,1579.1,301.00,666.52,761.65,0.0000,-3509.3,-6564.2,-290.52,-2616.3,-2450.8,-13601.,-1701.6,-1307.3,-5169.8,-2723.5,-5699.6,0.11173E+06,49943.,38258.,35906.,69606.,23986.,85976.,24845.,37982.,11337.,16293.,19626.,0.0000,-111.38,-115.74,-18.089,-106.50,-66.330,-436.15,-352.40,-36.177,-317.25,-38.205,-427.15
1604.000000000,8811.1,1613.0,1791.7,1637.0,2378.0,1125.5,2834.6,384.64,1567.2,302.35,673.36,762.63,0.0000,-3480.6,-6557.8,-288.53,-2616.7,-2430.9,-13601.,-1694.8,-1295.8,-5159.2,-2721.6,-5692.9,1296.9,579.68,444.05,416.76,807.90,278.40,997.91,288.37,440.85,131.59,189.12,227.80,0.0000,-1.2935,-1.3441,-0.20995,-1.2367,-0.77007,-5.0644,-4.0911,-0.41991,-3.6827,-0.44348,-4.9592
1605.000000000,8836.9,1651.3,1817.5,1626.6,2388.6,1157.3,2881.2,391.95,1559.9,306.17,691.89,776.49,0.0000,-3517.7,-6574.0,-290.37,-2617.4,-2456.3,-13604.,-1690.0,-1308.6,-5167.0,-2724.3,-5697.2,4021.1,1797.4,1376.8,1292.2,2505.0,863.20,3094.1,894.12,1366.9,408.00,586.37,706.31,0.0000,-4.0220,-4.1720,-0.65098,-3.8411,-2.4008,-15.715,-12.690,-1.3020,-11.421,-1.3757,-15.386
1606.000000000,8846.6,1606.2,1808.3,1627.0,2380.7,1117.1,2850.2,389.79,1537.0,305.25,691.41,776.19,0.0000,-3491.5,-6567.9,-288.52,-2617.5,-2437.1,-13605.,-1685.9,-1298.1,-5158.1,-2722.8,-5689.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1607.000000000,8934.6,1590.0,1788.0,1640.4,2381.4,1087.2,2799.2,387.73,1549.2,303.17,696.40,781.01,0.0000,-3483.1,-6556.8,-286.55,-2617.8,-2431.8,-13604.,-1682.9,-1292.6,-5154.2,-2722.8,-5684.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1608.000000000,9089.9,1582.9,1783.9,1644.9,2363.1,1068.1,2817.2,386.62,1546.2,300.14,701.13,785.47,0.0000,-3476.8,-6545.4,-284.99,-2618.0,-2428.3,-13602.,-1680.7,-1288.6,-5151.6,-2722.2,-5682.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1609.000000000,9084.2,1588.3,1795.7,1661.2,2353.6,1049.1,2819.5,376.43,1572.6,300.94,704.11,787.14,0.0000,-3471.5,-6535.6,-283.80,-2617.5,-2425.6,-13602.,-1679.2,-1285.5,-5149.7,-2721.9,-5680.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1610.000000000,9082.0,1577.9,1807.0,1684.4,2353.5,1066.0,2830.6,374.99,1581.7,298.46,704.84,783.22,0.0000,-3509.2,-6552.2,-286.90,-2616.6,-2450.1,-13602.,-1696.4,-1300.7,-5163.8,-2724.3,-5692.0,0.13595E+06,60767.,46549.,43688.,84691.,29184.,0.10461E+06,30229.,46214.,13794.,19825.,23880.,0.0000,-135.84,-140.98,-22.009,-129.77,-80.993,-531.09,-429.18,-44.018,-386.22,-46.492,-520.41
1611.000000000,9076.9,1593.2,1817.5,1691.4,2360.9,1068.3,2812.4,376.90,1582.5,300.34,703.47,781.72,0.0000,-3526.3,-6569.9,-290.04,-2616.0,-2458.6,-13601.,-1691.5,-1311.4,-5168.2,-2724.9,-5695.9,2421.8,1082.5,829.22,778.25,1508.7,519.88,1863.5,538.50,823.24,245.73,353.15,425.39,0.0000,-2.4237,-2.5130,-0.39206,-2.3132,-1.4441,-9.4598,-7.6457,-0.78413,-6.8800,-0.82821,-9.2702
1612.000000000,9120.1,1618.2,1818.1,1691.5,2374.9,1080.4,2864.8,381.45,1582.4,305.62,708.84,796.33,0.0000,-3540.5,-6587.0,-292.59,-2615.9,-2466.0,-13602.,-1746.8,-1319.8,-5181.1,-2725.8,-5712.3,0.44371E+06,0.19833E+06,0.15193E+06,0.14259E+06,0.27641E+06,95251.,0.34142E+06,98663.,0.15083E+06,45022.,64704.,77939.,0.0000,-444.99,-460.96,-71.833,-424.27,-265.02,-1734.1,-1401.9,-143.67,-1260.7,-151.74,-1699.2
1613.000000000,9131.0,1952.3,2024.5,1683.1,2510.8,1343.3,3205.7,419.14,1586.4,376.79,838.07,931.93,0.0000,-3570.2,-6616.8,-294.88,-2621.6,-2486.4,-13619.,-1735.3,-1327.1,-5197.4,-2737.6,-5721.3,51342.,22949.,17579.,16499.,31984.,11021.,39506.,11416.,17453.,5209.4,7486.8,9018.2,0.0000,-51.996,-53.527,-8.3117,-49.394,-31.292,-201.54,-162.54,-16.623,-146.07,-17.615,-197.23
1614.000000000,9171.4,1955.8,1973.6,1677.6,2509.4,1148.4,2946.9,409.26,1656.5,363.56,891.76,943.42,0.0000,-3590.3,-6637.1,-296.95,-2625.1,-2492.2,-13625.,-1720.5,-1334.4,-5202.4,-2749.9,-5723.7,10752.,4806.1,3681.6,3455.3,6698.3,2308.2,8273.7,2390.9,3655.1,1091.0,1568.0,1888.7,0.0000,-10.908,-11.215,-1.7407,-10.352,-6.5602,-42.202,-34.058,-3.4814,-30.598,-3.6893,-41.335
1615.000000000,9247.4,1970.9,1959.7,1659.2,2555.8,1104.0,2936.5,440.60,1688.3,350.76,927.58,925.20,0.0000,-3606.1,-6656.1,-298.78,-2625.2,-2496.6,-13629.,-1712.1,-1341.3,-5200.1,-2760.3,-5723.0,30562.,13661.,10465.,9821.3,19039.,6560.7,23517.,6795.7,10389.,3101.0,4456.7,5368.3,0.0000,-31.035,-31.894,-4.9478,-29.434,-18.631,-119.91,-96.832,-9.8955,-86.980,-10.486,-117.53
1616.000000000,9247.6,1915.9,1931.9,1642.5,2555.7,1106.3,3103.0,463.26,1712.0,351.73,857.16,879.58,0.0000,-3622.1,-6666.7,-300.38,-2624.2,-2500.3,-13634.,-1712.2,-1347.5,-5198.4,-2761.4,-5722.6,76671.,34270.,26252.,24638.,47763.,16459.,58996.,17048.,26063.,7779.4,11180.,13467.,0.0000,-77.972,-80.077,-12.412,-73.872,-46.709,-300.72,-242.98,-24.825,-218.23,-26.307,-294.90
1617.000000000,9254.8,1897.3,1933.7,1631.7,2579.9,1116.4,3107.4,453.60,1681.2,359.48,804.54,855.56,0.0000,-3636.6,-6676.6,-301.76,-2623.3,-2503.3,-13637.,-1703.7,-1353.0,-5196.5,-2758.9,-5721.6,10006.,4472.4,3426.0,3215.4,6233.1,2147.9,7699.1,2224.8,3401.3,1015.2,1459.1,1757.5,0.0000,-10.191,-10.459,-1.6198,-9.6436,-6.0910,-39.230,-31.713,-3.2397,-28.480,-3.4320,-38.488
1618.000000000,9193.0,1841.9,1976.4,1619.7,2649.9,1120.7,3072.2,443.31,1659.4,371.74,779.27,873.26,0.0000,-3604.8,-6662.8,-298.99,-2623.3,-2479.9,-13639.,-1696.1,-1335.4,-5182.5,-2753.3,-5712.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1619.000000000,9083.2,1822.9,1977.7,1621.4,2696.5,1106.4,2990.3,431.42,1645.1,365.16,818.71,879.53,0.0000,-3593.3,-6648.6,-296.31,-2623.6,-2473.6,-13641.,-1690.7,-1326.2,-5176.8,-2753.0,-5707.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1620.000000000,9044.9,1781.6,1986.6,1603.2,2617.4,1082.2,3012.0,428.89,1644.2,366.23,805.29,883.35,0.0000,-3584.3,-6636.9,-294.24,-2624.1,-2468.8,-13642.,-1686.8,-1320.6,-5174.6,-2753.5,-5704.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1621.000000000,9089.7,1791.5,1992.3,1600.3,2585.2,1063.6,3011.8,428.72,1655.0,359.03,786.32,873.50,0.0000,-3578.6,-6624.0,-292.69,-2624.7,-2464.5,-13643.,-1684.2,-1316.6,-5172.8,-2752.0,-5702.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1622.000000000,9133.0,1778.2,1970.4,1593.1,2680.1,1053.7,2983.5,421.17,1647.2,368.33,796.77,856.35,0.0000,-3571.8,-6612.6,-291.52,-2626.6,-2461.1,-13644.,-1682.3,-1312.3,-5172.5,-2750.9,-5700.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1623.000000000,9317.6,1809.9,1950.3,1607.6,2663.4,1069.0,2961.3,416.59,1660.6,363.05,797.72,849.65,0.0000,-3566.3,-6604.5,-290.64,-2628.1,-2458.1,-13644.,-1681.0,-1308.6,-5170.6,-2749.9,-5698.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1624.000000000,9490.6,1816.5,1931.0,1613.6,2636.7,1068.6,2981.8,413.52,1643.3,360.19,787.68,837.41,0.0000,-3561.7,-6597.2,-289.99,-2629.6,-2455.2,-13645.,-1680.1,-1305.3,-5168.9,-2748.5,-5696.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1625.000000000,9541.0,1791.9,1917.2,1617.9,2614.7,1090.7,3000.9,412.12,1650.5,361.49,783.20,830.28,0.0000,-3557.3,-6590.0,-289.47,-2632.0,-2453.4,-13645.,-1679.4,-1302.3,-5167.4,-2747.0,-5695.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1626.000000000,9554.7,1779.2,1890.4,1600.2,2601.0,1106.2,2992.7,405.46,1660.6,360.89,776.17,831.38,0.0000,-3553.1,-6583.4,-289.03,-2634.1,-2451.4,-13646.,-1678.9,-1299.5,-5166.2,-2746.0,-5694.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1627.000000000,9462.9,1764.1,1899.5,1614.7,2604.2,1103.5,3016.0,407.01,1647.7,361.07,773.24,828.65,0.0000,-3548.8,-6577.1,-288.64,-2635.5,-2449.2,-13646.,-1678.6,-1296.9,-5164.9,-2744.7,-5693.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1628.000000000,9435.6,1743.3,1892.7,1629.8,2620.6,1098.7,3015.6,419.05,1635.2,359.36,782.72,832.41,0.0000,-3544.1,-6570.6,-288.30,-2636.6,-2447.0,-13647.,-1678.4,-1294.5,-5163.5,-2744.0,-5692.8,694.91,310.61,237.94,223.31,432.90,149.18,534.71,154.52,236.22,70.509,101.33,122.06,0.0000,-0.70145,-0.72576,-0.11250,-0.66744,-0.41939,-2.7215,-2.2017,-0.22500,-1.9780,-0.23782,-2.6715
1629.000000000,9454.3,1753.5,1888.8,1649.4,2604.7,1104.5,3005.9,422.19,1621.6,360.27,780.46,846.67,0.0000,-3539.5,-6565.0,-287.98,-2637.6,-2444.8,-13647.,-1678.2,-1292.7,-5162.7,-2743.3,-5692.4,3.1112,1.3907,1.0653,0.99980,1.9382,0.66788,2.3940,0.69180,1.0576,0.31568,0.45369,0.54649,0.0000,-0.31383E-02,-0.32485E-02,-0.50368E-03,-0.29876E-02,-0.18771E-02,-0.12184E-01,-0.98562E-02,-0.10074E-02,-0.88551E-02,-0.10646E-02,-0.11959E-01
1630.000000000,9459.8,1725.7,1864.1,1653.8,2596.5,1091.2,3029.1,417.78,1626.8,358.79,777.75,857.65,0.0000,-3535.4,-6559.4,-287.67,-2638.4,-2442.7,-13648.,-1678.1,-1291.0,-5162.0,-2742.1,-5691.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1631.000000000,9469.1,1694.9,1854.7,1651.2,2594.2,1100.3,3035.7,416.61,1653.6,357.88,783.35,852.10,0.0000,-3531.2,-6554.5,-287.37,-2639.4,-2440.6,-13648.,-1677.9,-1289.4,-5161.3,-2740.8,-5691.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1632.000000000,9511.1,1663.1,1868.1,1651.9,2492.6,1115.2,3040.3,424.12,1670.7,359.23,783.16,846.68,0.0000,-3527.0,-6553.0,-287.08,-2640.4,-2438.5,-13648.,-1677.8,-1287.9,-5160.5,-2739.6,-5690.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1633.000000000,9639.0,1641.7,1835.0,1671.5,2449.6,1107.5,3054.2,424.42,1662.5,356.20,788.89,843.31,0.0000,-3523.0,-6551.2,-286.80,-2641.2,-2436.6,-13649.,-1677.7,-1286.5,-5159.7,-2738.6,-5690.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1634.000000000,9647.5,1621.9,1801.5,1673.2,2471.5,1122.6,3036.6,432.90,1645.5,356.63,783.81,849.47,0.0000,-3519.0,-6548.6,-286.53,-2641.9,-2434.8,-13649.,-1677.7,-1285.2,-5159.5,-2737.6,-5690.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1635.000000000,9560.0,1612.6,1791.4,1676.1,2471.4,1112.7,3028.0,426.85,1644.4,356.01,785.05,852.41,0.0000,-3515.0,-6545.4,-286.26,-2642.3,-2432.8,-13649.,-1677.6,-1283.9,-5159.1,-2736.6,-5689.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1636.000000000,9533.7,1615.6,1795.9,1671.1,2472.1,1115.5,3028.8,415.54,1641.3,355.38,782.92,846.76,0.0000,-3554.4,-6565.2,-289.98,-2642.7,-2458.1,-13650.,-1677.8,-1298.9,-5170.1,-2738.1,-5697.2,1685.9,753.57,577.25,541.77,1050.2,361.91,1297.2,374.87,573.09,171.06,245.84,296.13,0.0000,-1.6962,-1.7580,-0.27293,-1.6186,-1.0182,-6.5986,-5.3368,-0.54586,-4.7967,-0.57673,-6.4726
1637.000000000,9531.5,1591.5,1814.6,1677.2,2464.6,1119.1,2977.8,422.60,1645.0,356.04,766.23,840.37,0.0000,-3529.0,-6563.8,-289.56,-2643.2,-2439.5,-13649.,-1677.7,-1292.3,-5161.6,-2735.9,-5691.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1638.000000000,9482.9,1572.3,1810.4,1670.6,2428.3,1119.8,2984.7,427.10,1675.2,355.00,756.51,847.77,0.0000,-3521.4,-6559.5,-288.61,-2643.5,-2435.4,-13649.,-1677.8,-1288.9,-5158.7,-2734.7,-5689.8,1038.4,464.16,355.56,333.71,646.90,222.92,799.05,230.90,353.00,105.37,151.43,182.40,0.0000,-1.0438,-1.0828,-0.16811,-0.99682,-0.62628,-4.0636,-3.2865,-0.33623,-2.9543,-0.35520,-3.9855
1639.000000000,9467.4,1566.8,1815.9,1693.3,2418.3,1129.1,2989.2,428.83,1693.9,353.44,745.98,853.10,0.0000,-3559.3,-6577.6,-291.75,-2643.8,-2460.3,-13649.,-1682.7,-1303.6,-5169.7,-2736.4,-5698.4,37203.,16629.,12738.,11955.,23176.,7986.2,28626.,8272.3,12646.,3774.8,5425.0,6534.7,0.0000,-37.445,-38.810,-6.0228,-35.736,-22.488,-145.56,-117.73,-12.046,-105.84,-12.726,-142.76
1640.000000000,9483.3,1558.2,1802.5,1709.7,2404.0,1117.4,2988.6,424.42,1721.2,353.26,741.42,857.07,0.0000,-3576.6,-6596.0,-294.88,-2644.1,-2469.1,-13650.,-1682.4,-1314.5,-5173.1,-2736.8,-5702.0,7325.0,3274.1,2508.1,2353.9,4563.2,1572.4,5636.4,1628.8,2490.0,743.23,1068.2,1286.7,0.0000,-7.3844,-7.6470,-1.1859,-7.0417,-4.4353,-28.658,-23.179,-2.3717,-20.838,-2.5058,-28.105
1641.000000000,9486.8,1543.8,1766.4,1699.9,2395.0,1102.1,3020.2,419.86,1723.4,351.75,731.59,854.31,0.0000,-3546.7,-6589.8,-293.47,-2644.0,-2447.8,-13651.,-1681.0,-1304.2,-5162.4,-2734.3,-5695.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1642.000000000,9473.1,1540.6,1786.6,1715.2,2383.9,1091.5,3022.1,423.31,1715.9,352.01,731.59,851.72,0.0000,-3536.9,-6580.5,-291.72,-2643.9,-2442.3,-13653.,-1679.9,-1299.1,-5158.7,-2732.9,-5693.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1643.000000000,9450.0,1543.7,1786.7,1730.1,2352.8,1088.1,2993.2,422.89,1736.3,352.55,728.86,849.14,0.0000,-3530.0,-6571.8,-290.31,-2643.6,-2438.9,-13654.,-1679.1,-1296.1,-5156.8,-2731.6,-5691.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1644.000000000,9299.4,1578.6,1779.0,1735.7,2335.9,1093.4,2989.5,420.67,1756.1,350.15,722.92,840.77,0.0000,-3524.1,-6563.9,-289.23,-2643.3,-2436.0,-13655.,-1678.6,-1293.9,-5155.2,-2730.5,-5691.0,280.13,125.21,95.918,90.022,174.51,60.136,215.55,62.290,95.226,28.424,40.850,49.206,0.0000,-0.28181,-0.29234,-0.45351E-01,-0.26905,-0.16902,-1.0955,-0.88612,-0.90702E-01,-0.79676,-0.95798E-01,-1.0742
1645.000000000,9252.5,1550.2,1749.7,1744.0,2330.4,1118.3,2972.2,419.42,1746.3,346.96,722.69,832.70,0.0000,-3518.7,-6556.9,-288.39,-2643.0,-2433.4,-13655.,-1678.1,-1291.8,-5154.1,-2729.5,-5690.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1646.000000000,9196.3,1530.0,1744.9,1742.8,2321.6,1146.3,2948.7,420.25,1755.0,346.12,724.62,835.75,0.0000,-3513.5,-6550.8,-287.72,-2642.6,-2430.9,-13654.,-1677.8,-1290.0,-5153.1,-2728.7,-5689.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1647.000000000,9150.2,1574.7,1750.2,1748.6,2317.5,1171.3,2921.7,413.32,1794.7,348.87,714.56,841.60,0.0000,-3551.8,-6568.5,-291.16,-2642.2,-2456.0,-13653.,-1678.2,-1305.4,-5163.8,-2730.5,-5697.1,4370.4,1953.5,1496.4,1404.4,2722.6,938.18,3362.9,971.79,1485.6,443.44,637.31,767.67,0.0000,-4.3963,-4.5589,-0.70753,-4.1967,-2.6394,-17.084,-13.820,-1.4151,-12.429,-1.4944,-16.752
1648.000000000,9056.0,1586.7,1747.1,1761.9,2304.3,1193.5,2875.7,408.05,1814.9,349.85,707.11,844.15,0.0000,-3569.2,-6587.7,-294.51,-2641.9,-2464.6,-13653.,-1678.7,-1316.6,-5166.6,-2731.0,-5699.9,5667.0,2533.1,1940.4,1821.1,3530.3,1216.5,4360.6,1260.1,1926.4,575.01,826.39,995.43,0.0000,-5.7094,-5.9148,-0.91744,-5.4453,-3.4274,-22.150,-17.919,-1.8349,-16.116,-1.9378,-21.719
1649.000000000,9056.5,1568.3,1757.8,1786.8,2278.0,1184.3,2851.4,404.45,1798.4,346.82,699.87,845.93,0.0000,-3583.2,-6605.6,-297.20,-2641.5,-2471.1,-13652.,-1685.3,-1325.6,-5168.9,-2731.2,-5702.9,51924.,23209.,17779.,16686.,32346.,11146.,39954.,11546.,17651.,5268.5,7571.7,9120.6,0.0000,-52.402,-54.233,-8.4060,-49.927,-31.439,-202.92,-164.18,-16.812,-147.65,-17.755,-198.97
1650.000000000,9092.7,1568.7,1747.0,1794.8,2250.7,1181.3,2825.9,402.77,1792.7,342.28,692.75,836.49,0.0000,-3595.9,-6621.7,-299.32,-2641.2,-2476.8,-13651.,-1691.9,-1333.4,-5171.4,-2731.1,-5706.5,65017.,29061.,22262.,20893.,40502.,13957.,50028.,14457.,22101.,6596.9,9480.9,11420.,0.0000,-65.750,-67.961,-10.526,-62.560,-39.403,-254.05,-205.58,-21.051,-184.88,-22.231,-249.11
1651.000000000,9218.9,1558.4,1737.5,1780.7,2244.8,1158.1,2820.7,403.08,1776.8,342.71,691.93,833.20,0.0000,-3563.4,-6612.3,-297.03,-2640.9,-2454.3,-13649.,-1688.0,-1319.5,-5160.6,-2728.4,-5699.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1652.000000000,9213.9,1549.5,1722.2,1776.6,2253.1,1145.9,2824.0,404.02,1771.3,341.34,692.09,833.22,0.0000,-3551.5,-6599.6,-294.64,-2641.1,-2448.3,-13647.,-1684.9,-1312.5,-5156.6,-2727.0,-5696.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1653.000000000,9081.8,1549.7,1729.7,1782.1,2460.1,1157.4,2826.3,401.99,1768.3,337.85,691.56,832.72,0.0000,-3542.8,-6587.7,-292.76,-2641.3,-2444.9,-13646.,-1682.6,-1307.8,-5154.1,-2726.1,-5694.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1654.000000000,8924.4,1565.8,1794.9,1790.3,2477.0,1157.4,2828.0,402.51,1749.1,335.15,695.62,828.25,0.0000,-3536.3,-6577.3,-291.31,-2641.5,-2442.5,-13645.,-1680.9,-1304.1,-5152.3,-2725.4,-5692.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1655.000000000,8896.3,1558.6,1847.8,1805.2,2465.5,1157.8,2823.6,397.64,1731.1,332.02,703.27,820.04,0.0000,-3530.2,-6569.5,-290.17,-2641.3,-2439.6,-13644.,-1679.8,-1300.9,-5150.8,-2724.5,-5691.3,739.06,330.35,253.05,237.50,460.40,158.65,568.68,164.34,251.23,74.989,107.77,129.82,0.0000,-0.74518,-0.77205,-0.11965,-0.71037,-0.44647,-2.8879,-2.3367,-0.23929,-2.1015,-0.25265,-2.8315
1656.000000000,8885.0,1552.2,1847.2,1814.1,2452.2,1187.4,2811.4,400.21,1727.8,327.76,696.50,815.29,0.0000,-3567.9,-6585.0,-293.24,-2641.2,-2464.8,-13644.,-1680.4,-1316.9,-5161.6,-2726.3,-5698.2,10914.,4878.2,3736.8,3507.2,6798.8,2342.8,8397.7,2426.7,3709.9,1107.4,1591.5,1917.0,0.0000,-11.017,-11.404,-1.7668,-10.495,-6.6077,-42.642,-34.505,-3.5337,-31.033,-3.7309,-41.812
1657.000000000,8879.8,1543.6,1829.6,1831.2,2445.2,1205.9,2866.0,396.53,1728.3,325.29,689.57,809.12,0.0000,-3584.8,-6602.9,-296.30,-2641.2,-2473.3,-13642.,-1682.7,-1327.8,-5165.2,-2726.8,-5700.8,23527.,10516.,8055.8,7560.6,14657.,5050.6,18104.,5231.5,7997.7,2387.2,3430.8,4132.6,0.0000,-23.791,-24.597,-3.8089,-22.639,-14.267,-91.920,-74.386,-7.6177,-66.900,-8.0431,-90.134
1658.000000000,8868.9,1545.1,1815.2,1845.2,2424.1,1207.7,2891.9,397.45,1722.4,321.92,695.30,810.90,0.0000,-3598.2,-6619.6,-298.74,-2641.2,-2479.3,-13640.,-1686.2,-1336.1,-5167.4,-2726.9,-5702.9,36856.,16474.,12619.,11844.,22959.,7911.7,28359.,8195.1,12528.,3739.6,5374.4,6473.8,0.0000,-37.339,-38.557,-5.9666,-35.485,-22.366,-143.98,-116.52,-11.933,-104.80,-12.599,-141.19
1659.000000000,8859.0,1542.1,1809.7,1858.8,2405.9,1193.7,2859.9,398.85,1716.5,321.39,695.89,815.87,0.0000,-3610.1,-6634.4,-300.64,-2641.5,-2484.5,-13639.,-1686.1,-1343.2,-5168.6,-2727.0,-5704.0,17355.,7757.4,5942.4,5577.1,10811.,3725.6,13354.,3859.0,5899.5,1760.9,2530.8,3048.5,0.0000,-17.613,-18.169,-2.8096,-16.719,-10.537,-67.791,-54.869,-5.6193,-49.348,-5.9326,-66.479
1660.000000000,8788.1,1541.2,1812.9,1876.3,2400.0,1194.8,2856.3,398.64,1710.7,325.03,698.42,827.51,0.0000,-3621.1,-6647.2,-302.15,-2641.7,-2489.3,-13637.,-1684.7,-1349.5,-5169.2,-2726.9,-5704.3,7765.9,3471.2,2659.0,2495.6,4837.8,1667.1,5975.6,1726.8,2639.9,787.97,1132.5,1364.1,0.0000,-7.8955,-8.1366,-1.2572,-7.4860,-4.7173,-30.332,-24.551,-2.5145,-22.081,-2.6546,-29.745
1661.000000000,8748.8,1535.6,1807.3,1873.8,2408.3,1220.7,2852.2,394.67,1715.9,324.72,700.55,825.85,0.0000,-3631.4,-6660.0,-303.40,-2641.9,-2494.0,-13635.,-1683.4,-1355.1,-5168.9,-2726.7,-5704.2,6371.5,2847.9,2181.6,2047.5,3969.2,1367.8,4902.7,1416.8,2165.9,646.49,929.12,1119.2,0.0000,-6.4895,-6.6811,-1.0315,-6.1462,-3.8720,-24.885,-20.142,-2.0630,-18.116,-2.1779,-24.402
1662.000000000,8750.2,1538.4,1782.0,1856.9,2400.3,1207.9,2821.2,395.59,1714.6,321.41,695.70,825.24,0.0000,-3596.6,-6648.5,-300.47,-2641.9,-2470.7,-13632.,-1681.5,-1337.7,-5156.7,-2724.0,-5695.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1663.000000000,8816.1,1551.6,1777.0,1870.2,2382.7,1210.5,2811.2,393.09,1701.9,320.56,696.55,828.76,0.0000,-3582.9,-6633.3,-297.62,-2641.6,-2464.4,-13630.,-1680.1,-1328.6,-5152.3,-2722.8,-5692.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1664.000000000,9009.2,1567.7,1784.0,1878.7,2390.1,1217.8,2807.8,391.81,1690.1,322.28,699.79,829.73,0.0000,-3572.9,-6619.7,-295.41,-2640.9,-2460.3,-13628.,-1679.1,-1322.2,-5150.1,-2721.9,-5689.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1665.000000000,9014.9,1566.8,1789.0,1882.6,2384.4,1213.8,2812.5,387.17,1683.0,318.79,705.31,830.41,0.0000,-3564.6,-6608.2,-293.75,-2640.0,-2457.0,-13626.,-1678.5,-1317.0,-5148.7,-2721.4,-5688.1,500.77,223.83,171.46,160.92,311.96,107.50,385.32,111.35,170.23,50.810,73.024,87.961,0.0000,-0.50810,-0.52482,-0.81070E-01,-0.48241,-0.30281,-1.9559,-1.5828,-0.16214,-1.4238,-0.17112,-1.9175
1666.000000000,9052.0,1567.8,1807.5,1866.9,2377.1,1226.8,2810.4,390.72,1683.3,318.43,704.15,824.36,0.0000,-3601.0,-6620.6,-296.47,-2639.2,-2481.8,-13625.,-1695.2,-1333.0,-5162.7,-2723.5,-5699.0,0.12943E+06,57853.,44317.,41593.,80629.,27784.,99592.,28780.,43997.,13133.,18874.,22735.,0.0000,-131.50,-135.67,-20.954,-124.73,-78.411,-505.51,-409.16,-41.907,-367.99,-44.231,-495.59
1667.000000000,9153.3,1541.5,1843.8,1835.5,2386.8,1206.4,2833.5,393.12,1659.4,315.86,704.33,827.78,0.0000,-3572.4,-6612.2,-295.27,-2638.4,-2462.2,-13623.,-1690.6,-1321.7,-5155.5,-2721.6,-5694.7,1017.5,454.78,348.38,326.96,633.83,218.42,782.90,226.24,345.86,103.24,148.37,178.72,0.0000,-1.0328,-1.0664,-0.16472,-0.98016,-0.61541,-3.9736,-3.2165,-0.32943,-2.8927,-0.34766,-3.8957
1668.000000000,9144.5,1539.3,1788.3,1828.0,2408.9,1197.6,2873.4,390.96,1647.0,316.90,701.94,834.27,0.0000,-3561.9,-6601.2,-293.70,-2637.8,-2457.5,-13622.,-1686.8,-1315.4,-5152.4,-2721.1,-5692.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1669.000000000,9157.3,1561.0,1784.7,1832.9,2423.0,1206.2,2902.3,392.56,1627.4,318.66,712.23,834.01,0.0000,-3555.7,-6591.0,-292.39,-2637.5,-2455.4,-13622.,-1683.8,-1310.8,-5150.3,-2721.3,-5689.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1670.000000000,9165.9,1544.8,1766.2,1816.9,2451.4,1191.0,2886.4,388.28,1612.0,318.80,715.91,822.84,0.0000,-3549.6,-6582.2,-291.33,-2636.7,-2452.3,-13621.,-1681.7,-1306.9,-5149.1,-2720.9,-5687.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1671.000000000,9150.4,1549.5,1751.5,1813.7,2456.9,1204.0,2872.7,392.95,1600.2,320.34,709.24,819.22,0.0000,-3543.7,-6573.1,-290.44,-2636.3,-2449.2,-13620.,-1680.1,-1303.5,-5147.8,-2720.7,-5686.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1672.000000000,9141.3,1557.9,1750.6,1825.2,2450.9,1204.1,2859.6,391.01,1594.4,322.71,713.22,823.44,0.0000,-3537.9,-6565.1,-289.70,-2635.5,-2446.1,-13619.,-1679.1,-1300.4,-5146.6,-2720.2,-5684.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1673.000000000,9135.9,1543.6,1742.7,1832.0,2317.7,1211.5,2858.1,391.68,1608.9,321.18,722.04,821.82,0.0000,-3575.8,-6582.1,-293.06,-2634.7,-2470.6,-13619.,-1680.4,-1316.7,-5157.6,-2722.7,-5691.5,15538.,6945.0,5320.1,4993.1,9679.3,3335.4,11956.,3454.9,5281.7,1576.5,2265.7,2729.2,0.0000,-15.723,-16.255,-2.5154,-14.949,-9.3901,-60.678,-49.126,-5.0308,-44.181,-5.3080,-59.507
1674.000000000,9151.5,1529.0,1716.6,1835.3,2318.1,1209.9,2844.8,394.67,1623.4,320.73,725.04,825.79,0.0000,-3592.8,-6600.4,-296.32,-2634.1,-2478.8,-13618.,-1680.4,-1327.7,-5160.7,-2723.8,-5693.5,7458.2,3333.7,2553.7,2396.7,4646.1,1601.0,5738.8,1658.4,2535.3,756.75,1087.6,1310.0,0.0000,-7.5605,-7.8061,-1.2074,-7.1795,-4.5109,-29.121,-23.580,-2.4148,-21.207,-2.5480,-28.561
1675.000000000,9271.0,1525.6,1719.5,1841.8,2202.8,1199.0,2840.5,393.01,1625.2,318.82,725.50,827.16,0.0000,-3606.2,-6618.0,-298.93,-2633.6,-2484.9,-13617.,-1682.4,-1336.3,-5161.9,-2725.0,-5694.6,22074.,9866.6,7558.1,7093.5,13751.,4738.6,16985.,4908.3,7503.6,2239.7,3218.9,3877.3,0.0000,-22.419,-23.118,-3.5736,-21.262,-13.359,-86.176,-69.786,-7.1471,-62.764,-7.5416,-84.524
1676.000000000,9409.9,1532.3,1704.3,1847.5,2190.1,1202.0,2827.1,391.41,1613.8,318.79,718.45,823.75,0.0000,-3618.4,-6634.0,-300.95,-2633.0,-2490.3,-13615.,-1684.3,-1343.3,-5163.1,-2725.8,-5695.8,25403.,11355.,8698.0,8163.3,15825.,5453.2,19547.,5648.5,8635.2,2577.5,3704.3,4462.1,0.0000,-25.848,-26.623,-4.1125,-24.485,-15.380,-99.159,-80.309,-8.2250,-72.228,-8.6791,-97.263
1677.000000000,9370.0,1521.6,1686.6,1844.3,2209.3,1183.3,2867.9,396.82,1594.0,316.29,715.00,812.41,0.0000,-3585.5,-6624.7,-298.57,-2632.2,-2467.4,-13613.,-1682.2,-1327.6,-5151.8,-2723.5,-5687.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1678.000000000,9362.3,1519.5,1695.7,1863.2,2195.3,1197.1,2894.3,391.99,1614.7,312.73,720.64,816.71,0.0000,-3617.6,-6635.4,-300.07,-2631.6,-2488.8,-13613.,-1680.9,-1340.6,-5159.2,-2725.1,-5692.6,2056.4,919.19,704.12,660.85,1281.1,441.45,1582.4,457.26,699.05,208.66,299.88,361.22,0.0000,-2.0941,-2.1565,-0.33292,-1.9827,-1.2436,-8.0253,-6.5006,-0.66584,-5.8468,-0.70251,-7.8722
1679.000000000,9325.7,1500.1,1700.8,1839.7,2187.2,1177.1,2909.4,396.24,1637.8,311.74,718.99,816.93,0.0000,-3587.3,-6625.4,-297.87,-2631.0,-2467.7,-13611.,-1679.6,-1326.7,-5149.1,-2722.7,-5685.5,13.105,5.8576,4.4871,4.2113,8.1637,2.8132,10.084,2.9139,4.4547,1.3297,1.9110,2.3019,0.0000,-0.13333E-01,-0.13742E-01,-0.21215E-02,-0.12631E-01,-0.79092E-02,-0.51137E-01,-0.41423E-01,-0.42431E-02,-0.37258E-01,-0.44763E-02,-0.50161E-01
1680.000000000,9232.5,1481.9,1708.0,1826.0,2195.9,1177.6,2930.4,401.47,1641.2,311.19,712.50,814.46,0.0000,-3575.5,-6612.6,-295.59,-2630.3,-2461.8,-13611.,-1678.6,-1319.0,-5145.4,-2721.3,-5682.5,2.4611,1.1001,0.84267,0.79088,1.5331,0.52831,1.8937,0.54724,0.83660,0.24971,0.35888,0.43229,0.0000,-0.25010E-02,-0.25802E-02,-0.39843E-03,-0.23710E-02,-0.14831E-02,-0.96027E-02,-0.77788E-02,-0.79685E-03,-0.69969E-02,-0.84054E-03,-0.94191E-02
1681.000000000,9227.5,1477.3,1718.0,1818.6,2210.3,1214.4,2936.1,397.38,1657.0,314.08,707.80,815.96,0.0000,-3610.9,-6624.0,-297.75,-2629.7,-2485.4,-13612.,-1679.0,-1334.2,-5155.4,-2722.6,-5689.0,7988.2,3570.6,2735.2,2567.0,4976.3,1714.8,6146.7,1776.2,2715.4,810.53,1164.9,1403.1,0.0000,-8.1286,-8.3770,-1.2932,-7.6985,-4.8212,-31.165,-25.247,-2.5864,-22.710,-2.7281,-30.570
1682.000000000,9132.8,1474.9,1772.7,1804.4,2204.9,1204.6,2929.7,403.78,1686.8,314.49,702.93,812.13,0.0000,-3626.1,-6638.1,-300.12,-2629.2,-2492.9,-13612.,-1700.6,-1343.4,-5162.6,-2722.2,-5696.5,0.16691E+06,74605.,57150.,53637.,0.10398E+06,35830.,0.12843E+06,37113.,56738.,16935.,24339.,29318.,0.0000,-170.12,-175.13,-27.021,-160.94,-100.82,-651.10,-527.59,-54.042,-474.51,-57.001,-638.71
1683.000000000,9083.1,1479.5,1836.2,1792.2,2171.0,1188.0,2959.0,404.07,1673.7,315.31,700.51,806.51,0.0000,-3593.7,-6628.7,-298.07,-2628.7,-2470.5,-13611.,-1694.4,-1328.3,-5154.0,-2719.1,-5691.6,55.972,25.018,19.165,17.987,34.868,12.015,43.069,12.446,19.027,5.6792,8.1620,9.8316,0.0000,-0.57003E-01,-0.58732E-01,-0.90614E-02,-0.53952E-01,-0.33746E-01,-0.21834,-0.17694,-0.18123E-01,-0.15912,-0.19112E-01,-0.21419
1684.000000000,9116.3,1526.3,1859.8,1790.0,2152.9,1235.3,3011.7,414.16,1677.8,320.02,709.11,822.96,0.0000,-3627.7,-6639.7,-299.85,-2629.0,-2494.5,-13613.,-1689.6,-1341.8,-5162.3,-2721.4,-5696.9,1603.4,716.67,548.99,515.25,998.83,344.19,1233.7,356.52,545.03,162.69,233.81,281.63,0.0000,-1.6373,-1.6838,-0.25957,-1.5475,-0.97107,-6.2587,-5.0698,-0.51914,-4.5590,-0.54767,-6.1381
1685.000000000,9125.4,1514.1,1878.6,1780.8,2291.6,1203.0,3009.7,407.76,1659.0,319.38,715.40,818.69,0.0000,-3598.5,-6632.0,-297.87,-2629.0,-2474.6,-13614.,-1685.8,-1328.1,-5153.0,-2719.6,-5689.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1686.000000000,9106.6,1514.8,1862.5,1772.9,2221.6,1177.9,2971.5,403.46,1678.1,317.52,709.46,820.10,0.0000,-3587.1,-6620.2,-295.75,-2628.6,-2468.4,-13614.,-1682.9,-1320.7,-5150.1,-2718.9,-5685.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1687.000000000,8992.7,1521.3,1845.6,1762.8,2215.4,1166.4,2942.1,403.99,1680.6,314.96,713.40,821.08,0.0000,-3578.5,-6607.5,-294.02,-2628.5,-2463.9,-13613.,-1680.9,-1315.3,-5147.8,-2719.1,-5683.2,25.941,11.595,8.8820,8.3361,16.160,5.5686,19.960,5.7681,8.8180,2.6321,3.7827,4.5565,0.0000,-0.26411E-01,-0.27222E-01,-0.41995E-02,-0.25009E-01,-0.15673E-01,-0.10125,-0.82037E-01,-0.83991E-02,-0.73769E-01,-0.88585E-02,-0.99339E-01
1688.000000000,8911.9,1514.8,1840.0,1758.5,2181.5,1164.1,2939.3,400.32,1721.7,313.13,717.09,825.25,0.0000,-3570.8,-6596.6,-292.66,-2628.0,-2460.5,-13612.,-1679.5,-1311.1,-5146.0,-2719.4,-5681.7,1.6223,0.72513,0.55547,0.52132,1.0106,0.34825,1.2483,0.36072,0.55146,0.16460,0.23657,0.28496,0.0000,-0.16497E-02,-0.17017E-02,-0.26263E-03,-0.15632E-02,-0.97930E-03,-0.63315E-02,-0.51304E-02,-0.52526E-03,-0.46134E-02,-0.55396E-03,-0.62124E-02
1689.000000000,8975.6,1508.6,1852.8,1744.0,2170.5,1183.1,2934.3,402.91,1728.4,312.65,729.76,821.60,0.0000,-3607.7,-6612.1,-295.61,-2627.4,-2485.3,-13613.,-1680.2,-1327.4,-5157.0,-2722.7,-5688.6,11921.,5328.7,4081.9,3831.0,7426.6,2559.2,9173.2,2650.8,4052.5,1209.6,1738.4,2094.0,0.0000,-12.140,-12.507,-1.9300,-11.492,-7.2107,-46.524,-37.701,-3.8600,-33.902,-4.0713,-45.651
1690.000000000,8971.9,1522.9,1855.2,1747.4,2167.7,1171.5,2911.8,412.43,1726.5,311.96,732.79,816.00,0.0000,-3623.8,-6629.3,-298.60,-2626.8,-2493.4,-13613.,-1679.9,-1338.2,-5160.0,-2724.6,-5690.6,5702.0,2548.7,1952.4,1832.4,3552.1,1224.0,4387.5,1267.9,1938.3,578.56,831.49,1001.6,0.0000,-5.8162,-5.9848,-0.92310,-5.4990,-3.4517,-22.249,-18.031,-1.8462,-16.215,-1.9474,-21.833
1691.000000000,8897.9,1510.0,1839.6,1724.6,2161.2,1144.7,2891.9,407.45,1710.8,309.10,732.30,811.96,0.0000,-3592.3,-6622.3,-296.99,-2626.2,-2471.0,-13612.,-1678.9,-1324.6,-5149.3,-2723.2,-5683.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1692.000000000,8846.2,1479.6,1824.2,1754.0,2159.4,1129.8,2910.1,405.85,1718.9,309.20,718.64,802.87,0.0000,-3581.1,-6610.2,-295.05,-2625.7,-2464.8,-13611.,-1678.1,-1317.7,-5145.6,-2721.8,-5680.5,393.35,175.82,134.68,126.40,245.04,84.439,302.67,87.463,133.71,39.911,57.359,69.092,0.0000,-0.40034,-0.41270,-0.63679E-01,-0.37899,-0.23709,-1.5343,-1.2436,-0.12736,-1.1185,-0.13430,-1.5057
1693.000000000,9002.3,1472.6,1819.9,1768.8,2146.2,1146.7,2932.2,409.87,1733.3,311.66,718.13,800.29,0.0000,-3572.9,-6599.0,-293.44,-2625.1,-2460.6,-13611.,-1677.5,-1312.8,-5143.8,-2720.4,-5679.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1694.000000000,9168.1,1464.5,1807.2,1776.6,2168.7,1148.1,2927.1,406.53,1738.9,312.13,718.83,801.33,0.0000,-3565.6,-6588.3,-292.17,-2624.8,-2457.1,-13610.,-1677.0,-1308.8,-5142.4,-2719.3,-5677.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1695.000000000,9149.8,1456.2,1802.3,1770.6,2178.2,1143.8,2946.2,407.19,1734.6,314.65,716.21,797.92,0.0000,-3559.1,-6579.3,-291.16,-2624.4,-2453.9,-13610.,-1676.6,-1305.2,-5141.3,-2718.4,-5676.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1696.000000000,9087.8,1444.7,1789.5,1764.9,2173.6,1147.0,2959.0,403.11,1740.2,319.21,717.17,793.22,0.0000,-3552.9,-6571.8,-290.34,-2623.8,-2451.0,-13609.,-1676.4,-1301.9,-5140.3,-2717.4,-5676.0,118.91,53.149,40.714,38.211,74.074,25.526,91.496,26.440,40.420,12.065,17.340,20.886,0.0000,-0.12045,-0.12452,-0.19250E-01,-0.11435,-0.71320E-01,-0.46361,-0.37581,-0.38500E-01,-0.33804,-0.40582E-01,-0.45492
1697.000000000,9097.1,1451.6,1781.8,1766.4,2177.8,1178.4,2959.8,400.21,1759.5,319.56,710.38,790.04,0.0000,-3590.9,-6588.6,-293.63,-2623.3,-2476.1,-13609.,-1681.7,-1318.2,-5152.1,-2719.2,-5684.6,40931.,18295.,14015.,13153.,25498.,8786.5,31495.,9101.3,13914.,4153.1,5968.7,7189.6,0.0000,-41.522,-42.869,-6.6263,-39.379,-24.596,-159.57,-129.36,-13.253,-116.36,-13.969,-156.57
1698.000000000,9101.9,1458.7,1665.8,1746.8,2243.3,1190.9,2958.2,398.87,1750.3,318.12,702.51,793.98,0.0000,-3608.0,-6607.5,-296.84,-2623.4,-2484.5,-13609.,-1686.9,-1329.0,-5156.5,-2719.7,-5689.3,50013.,22355.,17125.,16072.,31156.,10736.,38484.,11121.,17001.,5074.6,7293.1,8784.9,0.0000,-50.825,-52.405,-8.0967,-48.145,-30.092,-194.96,-158.06,-16.193,-142.18,-17.069,-191.30
1699.000000000,8994.4,1460.5,1666.4,1737.9,2222.1,1203.0,2934.9,400.89,1748.9,319.02,708.91,800.73,0.0000,-3621.7,-6624.9,-299.38,-2623.3,-2490.8,-13609.,-1684.8,-1337.5,-5158.0,-2719.9,-5691.1,6158.1,2752.6,2108.5,1978.9,3836.2,1321.9,4738.5,1369.3,2093.3,624.83,898.00,1081.7,0.0000,-6.2694,-6.4565,-0.99694,-5.9319,-3.7090,-24.004,-19.461,-1.9939,-17.506,-2.1017,-23.552
1700.000000000,9117.7,1438.6,1654.3,1741.8,2227.7,1205.3,2896.0,403.93,1757.3,316.07,706.56,809.66,0.0000,-3633.7,-6639.6,-301.35,-2623.3,-2496.3,-13609.,-1686.5,-1344.6,-5158.9,-2720.3,-5692.5,31358.,14017.,10737.,10077.,19535.,6731.6,24129.,6972.7,10660.,3181.8,4572.8,5508.1,0.0000,-31.982,-32.900,-5.0766,-30.226,-18.903,-122.23,-99.099,-10.153,-89.140,-10.702,-119.92
1701.000000000,9199.8,1410.2,1641.8,1742.4,2220.3,1199.3,2901.5,403.77,1749.7,316.46,699.72,811.35,0.0000,-3600.0,-6628.8,-298.90,-2623.3,-2473.5,-13607.,-1683.6,-1328.8,-5147.6,-2717.9,-5684.8,470.85,210.46,161.22,151.31,293.32,101.08,362.31,104.70,160.06,47.775,68.661,82.706,0.0000,-0.47985,-0.49406,-0.76227E-01,-0.45376,-0.28329,-1.8352,-1.4879,-0.15245,-1.3384,-0.16066,-1.8005
1702.000000000,9164.1,1417.2,1641.5,1751.9,2189.7,1198.9,2899.7,400.32,1746.4,317.01,700.08,813.04,0.0000,-3587.0,-6615.2,-296.37,-2623.2,-2467.2,-13607.,-1681.3,-1320.6,-5143.5,-2716.6,-5681.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1703.000000000,9049.9,1423.3,1652.0,1748.4,2071.4,1191.0,2910.4,400.16,1747.5,316.02,698.89,812.09,0.0000,-3577.7,-6602.0,-294.36,-2622.8,-2463.3,-13607.,-1679.6,-1315.1,-5141.4,-2715.5,-5679.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1704.000000000,9018.9,1452.5,1670.1,1748.9,2080.8,1176.0,2907.9,404.96,1727.8,312.19,696.36,814.42,0.0000,-3570.2,-6590.7,-292.82,-2622.4,-2459.8,-13607.,-1678.4,-1310.6,-5139.9,-2714.3,-5678.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1705.000000000,9015.9,1465.7,1682.2,1758.6,2072.6,1187.0,2912.3,402.02,1714.0,312.75,702.59,814.65,0.0000,-3563.1,-6581.1,-291.63,-2621.9,-2456.8,-13607.,-1677.5,-1306.8,-5139.2,-2713.4,-5676.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1706.000000000,9004.3,1455.5,1675.3,1768.6,2071.8,1184.2,2898.6,399.88,1708.1,311.54,698.66,816.94,0.0000,-3556.3,-6572.7,-290.66,-2621.6,-2453.8,-13608.,-1676.9,-1303.5,-5139.0,-2712.6,-5675.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1707.000000000,9050.6,1457.5,1678.1,1779.6,2045.6,1192.0,2885.1,398.74,1712.7,315.32,690.53,815.84,0.0000,-3549.7,-6564.9,-289.86,-2621.5,-2451.0,-13608.,-1676.4,-1300.5,-5138.7,-2711.8,-5674.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1708.000000000,9155.5,1477.0,1678.4,1792.1,2027.7,1211.8,2855.3,397.88,1730.3,315.83,689.64,813.11,0.0000,-3587.8,-6581.0,-293.15,-2621.6,-2476.1,-13608.,-1676.4,-1316.8,-5149.9,-2714.0,-5681.7,1951.4,872.23,668.15,627.09,1215.6,418.90,1501.5,433.91,663.34,198.00,284.56,342.76,0.0000,-1.9793,-2.0433,-0.31591,-1.8774,-1.1731,-7.6082,-6.1653,-0.63182,-5.5466,-0.66563,-7.4606
1709.000000000,9271.5,1460.9,1674.6,1785.6,2020.6,1193.2,2863.8,394.92,1703.3,315.08,693.78,809.88,0.0000,-3560.8,-6577.7,-292.35,-2621.7,-2456.6,-13607.,-1676.1,-1307.6,-5141.7,-2712.2,-5675.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1710.000000000,9285.3,1458.9,1676.9,1775.0,2106.0,1172.0,2866.8,394.91,1704.1,312.89,694.31,812.05,0.0000,-3551.4,-6570.9,-291.07,-2621.6,-2451.7,-13606.,-1675.9,-1302.7,-5139.1,-2711.2,-5673.5,845.50,377.92,289.50,271.70,526.71,181.50,650.58,188.00,287.41,85.789,123.29,148.51,0.0000,-0.85605,-0.88483,-0.13688,-0.81290,-0.50704,-3.2960,-2.6709,-0.27376,-2.4031,-0.28835,-3.2319
1711.000000000,9288.8,1462.0,1676.7,1769.3,2141.0,1172.9,2872.8,396.39,1708.3,311.82,700.84,810.18,0.0000,-3544.6,-6563.8,-289.93,-2621.6,-2448.6,-13604.,-1675.7,-1299.2,-5137.8,-2710.7,-5672.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1712.000000000,9285.7,1454.3,1792.8,1755.4,2164.3,1181.3,2893.4,400.32,1703.3,310.26,711.04,807.78,0.0000,-3538.2,-6557.2,-289.01,-2621.6,-2446.0,-13603.,-1675.5,-1296.3,-5137.3,-2710.5,-5671.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1713.000000000,9290.5,1434.8,1802.8,1753.2,2168.2,1175.2,2906.0,399.84,1699.8,309.30,711.47,813.35,0.0000,-3532.3,-6550.0,-288.25,-2621.6,-2443.4,-13602.,-1675.3,-1293.7,-5137.0,-2710.5,-5671.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1714.000000000,9231.8,1440.3,1796.0,1752.3,2161.8,1171.2,2902.5,400.34,1687.6,308.70,709.48,819.74,0.0000,-3526.8,-6543.7,-287.61,-2621.3,-2441.0,-13601.,-1675.2,-1291.4,-5136.6,-2710.3,-5670.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1715.000000000,9115.1,1440.0,1793.3,1746.4,2159.9,1163.4,2889.2,393.47,1688.8,307.47,707.50,815.80,0.0000,-3521.4,-6538.0,-287.05,-2620.9,-2438.6,-13600.,-1675.1,-1289.3,-5136.1,-2710.2,-5670.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1716.000000000,9062.1,1435.3,1787.4,1743.3,2140.7,1140.1,2897.2,392.14,1687.5,308.71,703.16,811.57,0.0000,-3516.3,-6533.3,-286.53,-2620.3,-2436.3,-13599.,-1675.0,-1287.4,-5135.6,-2710.3,-5669.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1717.000000000,8908.4,1430.1,1796.3,1740.6,2125.3,1141.4,2912.1,395.39,1680.3,309.59,695.51,803.96,0.0000,-3511.3,-6528.7,-286.05,-2619.7,-2434.1,-13598.,-1674.9,-1285.7,-5135.1,-2709.9,-5669.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1718.000000000,8918.8,1425.8,1803.2,1752.4,2117.9,1158.7,2941.0,400.22,1674.0,310.59,690.46,805.82,0.0000,-3506.8,-6524.1,-285.59,-2619.1,-2431.9,-13597.,-1674.8,-1284.2,-5134.8,-2709.2,-5668.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1719.000000000,8890.4,1407.4,1799.8,1754.1,2116.4,1155.5,2925.5,402.77,1678.0,309.72,688.44,808.22,0.0000,-3502.5,-6519.6,-285.14,-2618.6,-2429.7,-13596.,-1674.7,-1282.7,-5134.3,-2708.4,-5668.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1720.000000000,8755.6,1400.7,1786.3,1754.7,2105.7,1156.3,2906.6,396.92,1672.9,308.41,688.39,808.07,0.0000,-3498.2,-6515.0,-284.71,-2618.0,-2427.5,-13596.,-1674.7,-1281.4,-5133.8,-2707.7,-5667.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1721.000000000,8743.8,1402.1,1775.9,1771.7,2100.9,1163.3,2902.7,390.92,1680.4,306.98,688.03,805.57,0.0000,-3494.2,-6511.0,-284.29,-2617.5,-2425.4,-13595.,-1674.6,-1279.9,-5133.3,-2706.9,-5667.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1722.000000000,8768.1,1390.8,1787.1,1769.6,2117.4,1168.5,2907.7,390.23,1678.6,308.71,688.55,799.16,0.0000,-3490.0,-6507.9,-283.89,-2616.9,-2423.4,-13595.,-1674.5,-1278.5,-5132.8,-2706.1,-5666.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1723.000000000,8791.8,1404.7,1788.6,1761.9,2146.4,1176.4,2919.7,391.64,1685.4,308.98,689.58,799.66,0.0000,-3485.8,-6505.2,-283.50,-2616.3,-2421.5,-13596.,-1674.4,-1277.4,-5132.3,-2705.5,-5665.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1724.000000000,8837.6,1405.4,1801.0,1768.2,2159.3,1194.7,2895.1,392.55,1698.5,308.00,693.71,799.30,0.0000,-3524.9,-6525.5,-287.08,-2615.8,-2447.1,-13597.,-1674.8,-1292.5,-5143.3,-2707.3,-5673.4,3088.6,1380.6,1057.5,992.54,1924.1,663.03,2376.6,686.78,1049.9,313.39,450.39,542.52,0.0000,-3.0975,-3.2135,-0.50002,-2.9567,-1.8379,-12.032,-9.7453,-1.0000,-8.7738,-1.0527,-11.791
1725.000000000,8934.4,1395.4,1783.7,1760.9,2144.1,1186.5,2886.8,394.41,1705.8,309.45,696.81,802.69,0.0000,-3499.9,-6524.6,-286.55,-2615.2,-2428.4,-13595.,-1674.7,-1286.3,-5134.9,-2705.5,-5667.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1726.000000000,9010.3,1385.9,1763.0,1762.7,2120.0,1184.6,2888.2,395.06,1710.3,310.86,694.99,804.81,0.0000,-3492.4,-6520.1,-285.48,-2614.4,-2424.3,-13594.,-1674.5,-1283.3,-5132.5,-2704.6,-5665.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1727.000000000,9062.3,1396.2,1756.9,1766.8,2130.6,1192.5,2921.9,392.09,1710.7,310.35,690.52,807.43,0.0000,-3530.5,-6538.5,-288.49,-2613.7,-2449.3,-13594.,-1674.8,-1298.2,-5142.9,-2706.4,-5672.9,2483.3,1110.0,850.27,798.00,1547.0,533.07,1910.8,552.17,844.13,251.96,362.12,436.19,0.0000,-2.4910,-2.5833,-0.40202,-2.3773,-1.4775,-9.6714,-7.8332,-0.80403,-7.0535,-0.84628,-9.4786
1728.000000000,9080.2,1407.9,1735.8,1763.7,2136.2,1186.7,2947.1,390.89,1707.0,310.88,688.98,813.18,0.0000,-3504.3,-6535.4,-287.54,-2613.1,-2430.3,-13592.,-1674.6,-1290.7,-5134.5,-2704.5,-5667.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1729.000000000,9082.4,1428.0,1746.6,1768.4,2130.6,1210.6,2928.7,393.52,1722.2,312.64,688.63,817.53,0.0000,-3539.2,-6551.8,-290.16,-2612.6,-2453.6,-13592.,-1693.9,-1304.6,-5147.6,-2706.1,-5678.4,0.14567E+06,65111.,49877.,46811.,90745.,31270.,0.11209E+06,32390.,49517.,14780.,21242.,25587.,0.0000,-146.25,-151.58,-23.582,-139.50,-86.711,-567.25,-459.51,-47.165,-413.74,-49.640,-555.97
1730.000000000,9136.7,1434.0,1769.8,1752.7,2124.3,1203.8,2905.9,398.36,1736.9,313.72,688.52,818.92,0.0000,-3555.4,-6570.0,-292.81,-2612.3,-2461.9,-13592.,-1700.4,-1314.7,-5154.5,-2706.5,-5685.8,85964.,38424.,29434.,27625.,53552.,18454.,66147.,19115.,29222.,8722.4,12536.,15100.,0.0000,-86.443,-89.512,-13.917,-82.379,-51.239,-334.73,-271.20,-27.834,-244.16,-29.295,-328.10
1731.000000000,9184.9,1432.6,1775.4,1763.3,2126.2,1202.3,2938.0,404.63,1714.3,317.31,684.96,828.57,0.0000,-3568.5,-6586.8,-294.98,-2611.7,-2468.4,-13592.,-1732.7,-1323.0,-5164.9,-2706.7,-5698.6,0.29283E+06,0.13089E+06,0.10026E+06,94102.,0.18242E+06,62861.,0.22532E+06,65113.,99542.,29712.,42701.,51436.,0.0000,-294.99,-305.22,-47.406,-280.84,-174.74,-1140.6,-924.30,-94.813,-831.77,-99.791,-1118.0
1732.000000000,9207.7,1639.0,1906.0,1772.0,2217.0,1397.3,3238.8,433.78,1715.5,351.19,749.25,900.95,0.0000,-3591.1,-6609.6,-296.90,-2614.7,-2485.4,-13602.,-1756.2,-1330.3,-5180.4,-2712.1,-5713.7,0.28844E+06,0.12893E+06,98763.,92692.,0.17969E+06,61919.,0.22195E+06,64138.,98051.,29267.,42062.,50666.,0.0000,-293.06,-301.55,-46.696,-277.98,-174.94,-1127.6,-912.26,-93.393,-820.15,-98.504,-1103.1
1733.000000000,9224.2,1807.4,2011.5,1777.4,2273.3,1422.7,3259.2,428.02,1710.2,399.74,831.54,985.25,0.0000,-3617.5,-6633.8,-298.66,-2620.9,-2498.8,-13614.,-1751.6,-1336.9,-5198.3,-2724.1,-5723.2,0.12968E+06,57964.,44402.,41673.,80785.,27838.,99784.,28835.,44082.,13158.,18910.,22778.,0.0000,-132.67,-135.86,-20.994,-125.42,-79.615,-508.26,-410.81,-41.988,-369.07,-44.363,-497.16
1734.000000000,9240.5,1844.8,1981.5,1776.7,2312.3,1306.6,3169.1,432.25,1783.9,384.99,915.94,995.38,0.0000,-3636.3,-6654.0,-300.42,-2624.4,-2505.3,-13622.,-1735.8,-1343.9,-5203.1,-2738.7,-5725.5,40584.,18140.,13896.,13042.,25282.,8712.1,31228.,9024.2,13796.,4117.9,5918.1,7128.7,0.0000,-41.612,-42.548,-6.5702,-39.292,-24.981,-159.11,-128.67,-13.140,-115.55,-13.891,-155.77
1735.000000000,9375.0,1869.0,1973.2,1775.2,2335.7,1269.1,3155.1,459.59,1795.2,378.34,957.70,989.93,0.0000,-3652.5,-6673.6,-302.08,-2625.2,-2510.5,-13628.,-1720.4,-1350.7,-5201.4,-2751.3,-5723.6,14099.,6301.9,4827.4,4530.7,8782.9,3026.5,10849.,3135.0,4792.6,1430.5,2055.9,2476.5,0.0000,-14.479,-14.791,-2.2825,-13.659,-8.6828,-55.266,-44.719,-4.5649,-40.151,-4.8277,-54.151
1736.000000000,9389.2,1845.4,1918.0,1763.1,2336.7,1208.0,3268.3,478.59,1802.4,370.49,907.87,950.93,0.0000,-3622.9,-6660.6,-299.59,-2624.2,-2485.3,-13632.,-1707.3,-1334.3,-5184.3,-2752.7,-5711.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1737.000000000,9418.0,1859.7,1910.5,1757.3,2371.3,1210.1,3355.5,488.53,1797.3,386.37,849.23,927.68,0.0000,-3614.0,-6644.1,-297.13,-2622.5,-2477.1,-13636.,-1698.0,-1326.1,-5176.6,-2750.6,-5704.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1738.000000000,9406.6,1794.3,1977.3,1753.7,2399.6,1252.9,3293.8,468.21,1803.6,396.53,802.26,929.49,0.0000,-3652.0,-6652.7,-299.23,-2621.2,-2498.8,-13640.,-1703.0,-1341.9,-5185.5,-2748.8,-5711.8,84977.,37983.,29096.,27308.,52937.,18242.,65387.,18895.,28886.,8622.2,12392.,14926.,0.0000,-87.077,-89.170,-13.757,-82.188,-51.966,-332.65,-269.64,-27.514,-242.05,-29.074,-326.51
1739.000000000,9410.0,1735.9,2012.1,1752.9,2458.2,1246.6,3246.8,460.27,1795.7,388.18,817.57,942.38,0.0000,-3667.5,-6663.8,-301.59,-2620.7,-2505.0,-13642.,-1697.6,-1351.3,-5186.7,-2748.6,-5714.0,14005.,6260.2,4795.4,4500.7,8724.8,3006.5,10777.,3114.2,4760.9,1421.1,2042.3,2460.1,0.0000,-14.371,-14.708,-2.2674,-13.549,-8.5672,-54.806,-44.441,-4.5347,-39.894,-4.7898,-53.812
1740.000000000,9414.2,1667.8,2041.5,1745.5,2390.0,1246.1,3253.0,454.50,1807.8,385.16,798.66,946.41,0.0000,-3634.3,-6654.9,-299.56,-2620.7,-2481.7,-13643.,-1691.7,-1336.9,-5175.1,-2745.7,-5706.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1741.000000000,9412.8,1650.8,2075.0,1735.3,2373.6,1268.0,3259.5,455.48,1800.5,381.13,799.14,953.23,0.0000,-3624.0,-6642.6,-297.36,-2621.3,-2476.1,-13646.,-1687.4,-1330.2,-5171.6,-2744.0,-5702.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1742.000000000,9409.2,1627.7,2057.1,1729.2,2456.3,1274.1,3242.1,448.09,1775.8,387.46,798.33,931.29,0.0000,-3616.1,-6632.1,-295.59,-2623.8,-2472.3,-13648.,-1684.4,-1324.9,-5170.7,-2742.3,-5699.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1743.000000000,9437.9,1661.1,2054.2,1703.6,2424.2,1312.6,3212.9,444.26,1814.9,384.33,790.48,915.62,0.0000,-3609.9,-6623.7,-294.21,-2626.0,-2469.0,-13649.,-1682.2,-1320.4,-5168.4,-2740.4,-5696.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1744.000000000,9570.9,1661.8,2032.8,1712.7,2395.0,1321.7,3185.0,438.17,1802.8,381.08,774.96,901.44,0.0000,-3648.5,-6638.5,-297.10,-2629.0,-2494.0,-13651.,-1686.7,-1336.8,-5178.7,-2741.0,-5703.6,44704.,19982.,15307.,14366.,27848.,9596.4,34398.,9940.2,15196.,4535.9,6518.8,7852.3,0.0000,-45.793,-46.980,-7.2371,-43.202,-27.293,-174.94,-141.85,-14.474,-127.35,-15.271,-171.75
1745.000000000,9606.0,1637.1,2001.0,1727.1,2377.2,1369.0,3160.5,437.25,1802.0,385.76,767.44,903.81,0.0000,-3666.2,-6654.0,-300.04,-2632.2,-2503.8,-13653.,-1684.6,-1347.0,-5180.7,-2741.2,-5705.5,2510.4,1122.1,859.57,806.74,1563.9,538.91,1931.7,558.21,853.37,254.72,366.08,440.96,0.0000,-2.5763,-2.6399,-0.40642,-2.4276,-1.5350,-9.8233,-7.9653,-0.81283,-7.1513,-0.85754,-9.6439
1746.000000000,9610.4,1633.5,1996.9,1714.0,2356.6,1342.9,3125.8,448.39,1832.9,383.15,764.57,909.02,0.0000,-3634.9,-6644.7,-298.42,-2634.5,-2482.6,-13653.,-1682.5,-1332.6,-5169.0,-2739.0,-5697.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1747.000000000,9587.0,1640.5,1973.8,1708.6,2340.9,1326.6,3166.2,440.31,1818.1,377.86,770.31,898.38,0.0000,-3623.4,-6632.3,-296.49,-2636.0,-2477.0,-13654.,-1681.0,-1325.4,-5164.1,-2738.1,-5694.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1748.000000000,9626.0,1640.5,1947.1,1703.1,2370.8,1310.8,3180.2,431.66,1806.7,375.41,763.57,896.99,0.0000,-3614.9,-6619.4,-294.91,-2637.3,-2473.0,-13655.,-1679.8,-1320.6,-5161.3,-2737.1,-5692.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1749.000000000,9617.9,1649.0,1946.2,1710.9,2336.6,1287.9,3162.3,428.43,1811.1,371.98,771.06,898.02,0.0000,-3607.2,-6607.4,-293.66,-2638.2,-2469.4,-13656.,-1679.0,-1316.7,-5159.3,-2735.7,-5690.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1750.000000000,9615.5,1652.3,1922.6,1711.6,2331.4,1279.7,3149.7,427.72,1806.7,368.11,766.81,891.84,0.0000,-3600.2,-6596.8,-292.67,-2639.1,-2466.2,-13657.,-1678.5,-1313.5,-5157.6,-2734.2,-5689.7,793.75,354.79,271.78,255.07,494.47,170.39,610.76,176.50,269.82,80.538,115.75,139.42,0.0000,-0.81051,-0.83377,-0.12850,-0.76636,-0.48294,-3.1052,-2.5173,-0.25700,-2.2605,-0.27098,-3.0469
1751.000000000,9616.3,1621.6,1920.7,1722.9,2310.1,1287.4,3133.7,434.30,1793.6,373.42,767.86,889.80,0.0000,-3593.9,-6589.2,-291.85,-2639.9,-2463.4,-13658.,-1678.1,-1310.7,-5156.2,-2732.7,-5688.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1752.000000000,9597.1,1601.5,1943.1,1731.9,2333.6,1282.1,3149.0,435.39,1790.3,372.59,774.40,886.74,0.0000,-3587.9,-6584.5,-291.15,-2640.6,-2460.6,-13658.,-1677.7,-1308.1,-5155.1,-2731.3,-5687.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1753.000000000,9591.9,1602.0,1934.4,1759.3,2336.4,1281.5,3150.4,440.39,1763.4,368.38,789.28,885.12,0.0000,-3581.8,-6578.7,-290.54,-2641.0,-2457.8,-13658.,-1677.5,-1305.7,-5154.7,-2730.2,-5686.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1754.000000000,9600.2,1605.7,1919.3,1763.1,2338.1,1297.1,3136.4,434.95,1755.1,370.40,781.97,884.17,0.0000,-3575.7,-6572.7,-289.98,-2641.4,-2455.1,-13658.,-1677.3,-1303.6,-5154.3,-2729.2,-5686.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1755.000000000,9581.6,1590.7,1908.4,1764.8,2323.4,1302.1,3120.2,430.25,1773.4,369.14,780.46,877.70,0.0000,-3570.1,-6567.4,-289.47,-2641.6,-2452.4,-13658.,-1677.2,-1301.6,-5153.7,-2728.4,-5685.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1756.000000000,9544.1,1562.3,1913.8,1758.9,2306.8,1307.4,3139.7,429.50,1790.2,368.37,781.80,871.73,0.0000,-3564.6,-6562.9,-288.99,-2641.9,-2449.8,-13658.,-1677.1,-1299.8,-5153.3,-2727.7,-5685.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1757.000000000,9475.1,1536.9,1937.8,1761.3,2345.0,1311.7,3116.7,435.95,1812.4,367.33,780.02,874.98,0.0000,-3559.1,-6558.8,-288.54,-2642.1,-2447.3,-13658.,-1677.0,-1298.1,-5152.9,-2726.9,-5685.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1758.000000000,9450.2,1522.0,1956.8,1777.9,2327.0,1302.0,3113.8,445.46,1810.9,368.11,774.89,876.88,0.0000,-3553.8,-6554.9,-288.11,-2642.1,-2444.8,-13657.,-1676.9,-1296.5,-5152.5,-2726.1,-5684.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1759.000000000,9444.0,1508.4,1953.3,1776.3,2381.5,1273.7,3120.3,442.81,1806.3,364.72,768.37,877.00,0.0000,-3548.7,-6550.9,-287.69,-2642.0,-2442.5,-13656.,-1676.8,-1295.2,-5152.1,-2725.4,-5683.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1760.000000000,9427.1,1508.5,1938.4,1767.5,2414.7,1266.0,3115.6,439.58,1804.9,363.34,763.62,878.85,0.0000,-3543.8,-6547.1,-287.30,-2641.9,-2440.3,-13654.,-1676.8,-1294.1,-5151.6,-2724.6,-5683.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1761.000000000,9418.8,1488.2,1925.2,1760.9,2388.6,1275.9,3122.2,441.27,1815.1,363.07,761.67,873.42,0.0000,-3539.1,-6542.7,-286.91,-2641.7,-2438.2,-13653.,-1676.7,-1292.9,-5150.9,-2723.6,-5683.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1762.000000000,9377.1,1503.1,1907.1,1771.1,2373.4,1288.9,3164.8,444.86,1828.5,364.08,755.97,868.15,0.0000,-3534.6,-6538.5,-286.52,-2641.6,-2436.3,-13653.,-1676.7,-1291.6,-5150.1,-2722.8,-5682.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1763.000000000,9435.8,1501.3,1894.7,1756.2,2369.8,1294.1,3182.8,441.53,1836.9,360.69,760.88,858.53,0.0000,-3529.9,-6535.1,-286.14,-2641.3,-2434.4,-13654.,-1676.6,-1290.4,-5149.4,-2722.3,-5682.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1764.000000000,9407.9,1494.3,1875.7,1753.0,2363.7,1298.7,3198.4,438.80,1836.1,356.95,758.25,859.26,0.0000,-3525.4,-6531.6,-285.79,-2641.0,-2432.4,-13654.,-1676.6,-1289.5,-5148.5,-2721.7,-5681.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1765.000000000,9394.8,1483.1,1864.2,1762.2,2349.1,1298.5,3207.5,437.85,1813.7,356.08,754.74,862.31,0.0000,-3521.1,-6528.2,-285.46,-2640.4,-2430.4,-13653.,-1676.5,-1288.6,-5147.7,-2721.0,-5681.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1766.000000000,9379.5,1483.7,1852.1,1766.0,2341.6,1305.8,3196.5,437.58,1797.8,361.79,755.78,861.86,0.0000,-3516.5,-6524.8,-285.10,-2639.8,-2428.4,-13651.,-1676.6,-1287.7,-5147.0,-2720.4,-5681.1,762.52,340.83,261.09,245.04,475.02,163.69,586.74,169.55,259.21,77.370,111.19,133.94,0.0000,-0.76725,-0.79617,-0.12345,-0.73236,-0.46018,-2.9814,-2.4139,-0.24689,-2.1697,-0.26011,-2.9191
1767.000000000,9271.3,1493.3,1859.2,1765.1,2331.9,1314.4,3189.6,436.75,1797.8,364.89,758.84,860.17,0.0000,-3512.0,-6521.5,-284.73,-2639.1,-2426.4,-13650.,-1676.5,-1286.8,-5146.3,-2719.8,-5680.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1768.000000000,9306.8,1477.7,1859.8,1773.9,2313.2,1316.5,3189.9,437.02,1809.8,363.51,758.34,859.97,0.0000,-3507.7,-6518.6,-284.36,-2638.1,-2424.6,-13649.,-1676.4,-1286.0,-5145.8,-2719.2,-5680.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1769.000000000,9301.1,1476.5,1857.2,1774.4,2314.8,1312.6,3198.5,436.33,1816.3,361.20,752.33,856.97,0.0000,-3503.5,-6515.9,-283.99,-2637.5,-2422.5,-13647.,-1676.4,-1285.2,-5145.3,-2718.5,-5680.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1770.000000000,9299.7,1484.1,1851.9,1767.2,2323.6,1304.8,3206.2,436.27,1799.8,359.78,750.78,857.17,0.0000,-3499.4,-6513.5,-283.62,-2637.0,-2420.6,-13646.,-1676.3,-1284.4,-5144.9,-2717.8,-5679.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1771.000000000,9294.4,1482.3,1845.9,1772.0,2320.8,1306.3,3224.2,440.34,1795.1,361.49,751.16,858.38,0.0000,-3495.5,-6511.1,-283.25,-2636.5,-2418.8,-13644.,-1676.3,-1283.6,-5144.5,-2717.1,-5678.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1772.000000000,9290.6,1485.4,1852.8,1799.6,2308.3,1302.1,3249.5,435.89,1790.9,362.71,751.25,864.17,0.0000,-3491.6,-6509.0,-282.89,-2636.0,-2416.9,-13643.,-1676.2,-1282.8,-5144.1,-2716.5,-5678.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1773.000000000,9294.5,1490.3,1860.3,1833.3,2294.7,1307.2,3249.6,439.86,1795.7,361.53,755.41,866.78,0.0000,-3487.7,-6507.3,-282.52,-2635.4,-2415.1,-13641.,-1676.2,-1282.0,-5143.9,-2715.9,-5677.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1774.000000000,9340.8,1483.5,1877.1,1851.5,2302.0,1339.3,3236.8,440.03,1803.2,360.97,757.49,862.87,0.0000,-3526.8,-6529.3,-286.13,-2634.7,-2440.5,-13641.,-1676.4,-1296.9,-5155.0,-2717.9,-5685.5,1704.6,761.93,583.66,547.79,1061.9,365.93,1311.7,379.03,579.45,172.96,248.57,299.42,0.0000,-1.7091,-1.7754,-0.27596,-1.6339,-1.0264,-6.6626,-5.3916,-0.55193,-4.8485,-0.58126,-6.5204
1775.000000000,9398.6,1474.7,1879.5,1834.7,2295.9,1335.7,3242.6,436.43,1796.0,359.09,760.55,861.61,0.0000,-3501.7,-6530.1,-285.60,-2633.9,-2422.1,-13639.,-1676.3,-1291.1,-5146.8,-2716.0,-5680.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1776.000000000,9404.0,1473.9,1883.2,1845.0,2281.9,1339.9,3244.0,437.89,1796.2,357.20,755.73,862.99,0.0000,-3494.5,-6526.7,-284.55,-2633.0,-2418.4,-13637.,-1676.2,-1288.2,-5144.3,-2715.1,-5678.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1777.000000000,9396.1,1474.1,1886.3,1868.4,2260.7,1363.5,3240.7,441.83,1800.5,357.44,754.17,867.04,0.0000,-3532.5,-6545.4,-287.55,-2632.2,-2443.4,-13637.,-1677.9,-1303.0,-5154.9,-2717.0,-5685.6,13353.,5968.7,4572.2,4291.1,8318.5,2866.5,10275.,2969.2,4539.2,1354.9,1947.2,2345.5,0.0000,-13.394,-13.908,-2.1618,-12.799,-8.0368,-52.188,-42.223,-4.3235,-37.975,-4.5527,-51.066
1778.000000000,9378.6,1469.4,1874.8,1856.0,2256.1,1369.1,3257.9,441.71,1793.5,358.43,752.80,870.80,0.0000,-3506.5,-6543.0,-286.59,-2631.4,-2424.8,-13635.,-1677.4,-1296.0,-5146.4,-2715.0,-5680.2,0.59471E-01,0.26583E-01,0.20363E-01,0.19111E-01,0.37048E-01,0.12767E-01,0.45761E-01,0.13224E-01,0.20216E-01,0.60343E-02,0.86723E-02,0.10446E-01,0.0000,-0.59633E-04,-0.61942E-04,-0.96279E-05,-0.56986E-04,-0.35742E-04,-0.23242E-03,-0.18803E-03,-0.19256E-04,-0.16912E-03,-0.20275E-04,-0.22741E-03
1779.000000000,9370.9,1476.0,1875.0,1851.4,2258.5,1382.5,3266.8,443.43,1805.7,356.57,757.34,870.07,0.0000,-3541.8,-6560.4,-289.20,-2630.5,-2448.4,-13635.,-1677.5,-1310.1,-5155.1,-2716.4,-5686.3,3751.1,1676.7,1284.4,1205.4,2336.8,805.23,2886.3,834.08,1275.1,380.60,546.99,658.88,0.0000,-3.7665,-3.9086,-0.60727,-3.5962,-2.2580,-14.659,-11.859,-1.2145,-10.667,-1.2788,-14.343
1780.000000000,9372.3,1465.0,1862.5,1839.7,2256.9,1364.2,3255.0,442.63,1798.9,356.58,754.81,862.43,0.0000,-3514.7,-6556.2,-287.87,-2629.5,-2429.0,-13634.,-1677.1,-1301.6,-5145.7,-2714.0,-5680.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1781.000000000,9380.0,1463.5,1845.9,1829.7,2257.4,1360.5,3249.4,445.30,1788.8,357.16,751.00,855.94,0.0000,-3505.9,-6548.6,-286.25,-2628.5,-2424.4,-13632.,-1676.7,-1297.3,-5142.5,-2712.8,-5677.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1782.000000000,9375.0,1470.2,1820.5,1816.7,2253.6,1369.3,3251.2,443.65,1791.1,357.16,749.76,856.80,0.0000,-3499.5,-6541.3,-284.92,-2627.4,-2421.6,-13631.,-1676.3,-1294.3,-5141.1,-2711.8,-5676.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1783.000000000,9357.6,1481.4,1817.8,1825.7,2252.1,1359.9,3246.3,441.37,1789.1,358.15,750.11,852.87,0.0000,-3493.7,-6534.6,-283.87,-2626.4,-2419.1,-13630.,-1676.1,-1291.9,-5140.1,-2711.0,-5675.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1784.000000000,9339.1,1470.1,1843.5,1839.3,2254.2,1359.5,3232.8,440.67,1827.6,358.38,752.53,854.20,0.0000,-3488.4,-6529.1,-283.03,-2625.4,-2417.0,-13630.,-1675.9,-1289.9,-5139.4,-2710.3,-5675.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1785.000000000,9329.8,1467.5,1835.9,1846.8,2257.8,1363.7,3221.0,446.80,1857.3,355.40,757.91,853.49,0.0000,-3483.6,-6524.3,-282.35,-2624.5,-2414.9,-13629.,-1675.7,-1288.2,-5138.5,-2709.7,-5674.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1786.000000000,9338.8,1475.4,1829.0,1854.1,2193.9,1359.6,3201.3,445.19,1858.4,353.37,760.70,858.21,0.0000,-3479.0,-6520.0,-281.77,-2623.4,-2412.9,-13628.,-1675.6,-1286.6,-5137.7,-2709.1,-5673.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1787.000000000,9340.8,1453.5,1815.3,1863.3,2136.2,1345.4,3171.9,452.33,1855.3,354.66,760.43,859.64,0.0000,-3474.5,-6515.9,-281.26,-2622.3,-2410.8,-13626.,-1675.5,-1285.3,-5136.9,-2708.5,-5673.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1788.000000000,9358.9,1446.7,1800.8,1878.5,2119.6,1350.7,3176.2,451.78,1864.5,351.52,755.80,862.55,0.0000,-3470.1,-6512.2,-280.80,-2621.3,-2408.8,-13625.,-1675.4,-1283.9,-5136.4,-2708.0,-5672.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1789.000000000,9359.5,1448.7,1792.7,1875.6,2119.0,1354.8,3179.8,447.10,1860.9,347.89,757.64,868.61,0.0000,-3465.7,-6508.4,-280.42,-2620.3,-2406.8,-13624.,-1675.3,-1282.6,-5135.9,-2707.4,-5672.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1790.000000000,9375.7,1450.1,1797.7,1873.7,2125.8,1350.2,3194.6,448.49,1856.4,346.95,756.62,872.13,0.0000,-3461.4,-6504.9,-280.06,-2619.3,-2404.9,-13623.,-1675.2,-1281.4,-5135.4,-2706.9,-5672.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1791.000000000,9374.4,1441.7,1845.1,1864.0,2118.6,1341.2,3203.8,451.30,1853.5,347.09,756.30,875.78,0.0000,-3457.3,-6501.5,-279.71,-2618.3,-2403.0,-13622.,-1675.1,-1280.3,-5135.0,-2706.5,-5671.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1792.000000000,9369.3,1431.4,1900.7,1866.5,2123.0,1340.2,3194.3,453.19,1826.8,345.67,756.18,877.31,0.0000,-3453.3,-6498.2,-279.37,-2617.3,-2401.1,-13620.,-1675.1,-1279.2,-5134.5,-2706.0,-5671.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1793.000000000,9398.7,1425.9,1894.1,1873.4,2128.0,1327.4,3193.1,457.60,1828.5,344.55,752.34,872.89,0.0000,-3449.4,-6495.0,-279.05,-2616.2,-2399.2,-13619.,-1675.0,-1278.2,-5134.0,-2705.5,-5671.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1794.000000000,9408.9,1442.2,1888.9,1879.7,2131.6,1328.0,3199.0,460.50,1842.0,344.31,746.24,871.01,0.0000,-3445.6,-6492.0,-278.73,-2615.1,-2397.3,-13617.,-1674.9,-1277.3,-5133.4,-2705.0,-5670.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1795.000000000,9269.6,1457.8,1895.4,1872.1,2150.2,1324.4,3194.9,459.24,1816.5,341.77,744.75,868.73,0.0000,-3441.9,-6489.3,-278.43,-2614.0,-2395.5,-13616.,-1674.8,-1276.3,-5132.8,-2704.4,-5670.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1796.000000000,9116.1,1453.3,1902.3,1864.9,2154.1,1314.2,3171.8,460.31,1809.7,343.25,746.73,866.11,0.0000,-3438.2,-6486.6,-278.12,-2612.8,-2393.8,-13615.,-1674.8,-1275.4,-5132.3,-2703.9,-5670.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1797.000000000,9138.6,1443.2,1901.9,1852.6,2136.2,1319.2,3179.1,460.56,1803.1,345.03,749.23,861.89,0.0000,-3434.5,-6484.1,-277.81,-2611.7,-2392.1,-13614.,-1674.7,-1274.5,-5131.9,-2703.4,-5670.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1798.000000000,9129.9,1444.1,1886.4,1840.5,2145.2,1320.1,3179.4,461.12,1814.7,345.44,749.88,858.34,0.0000,-3430.9,-6481.7,-277.50,-2610.6,-2390.4,-13612.,-1674.6,-1273.7,-5131.4,-2702.9,-5669.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1799.000000000,9133.9,1443.4,1876.8,1832.3,2135.4,1301.6,3168.7,461.74,1836.8,347.82,747.78,853.32,0.0000,-3427.5,-6479.6,-277.19,-2609.5,-2388.7,-13611.,-1674.5,-1272.9,-5131.0,-2702.4,-5669.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1800.000000000,9113.6,1437.0,1870.1,1835.3,2130.8,1307.0,3178.1,460.72,1838.8,350.48,743.73,853.82,0.0000,-3424.0,-6477.7,-276.88,-2608.4,-2387.1,-13609.,-1674.5,-1272.2,-5130.6,-2701.8,-5669.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1801.000000000,9122.8,1421.4,1773.5,1836.0,2135.1,1335.8,3188.1,456.97,1840.9,352.07,744.74,850.91,0.0000,-3463.4,-6498.8,-280.53,-2607.4,-2412.8,-13608.,-1679.7,-1286.1,-5142.7,-2703.9,-5678.3,39033.,17447.,13365.,12543.,24316.,8379.1,30035.,8679.3,13269.,3960.5,5691.9,6856.2,0.0000,-38.731,-40.367,-6.3191,-37.169,-23.113,-152.39,-123.15,-12.638,-110.88,-13.290,-149.01
1802.000000000,9092.3,1441.5,1754.1,1848.9,2126.9,1328.8,3193.5,459.02,1854.8,353.74,745.92,854.03,0.0000,-3481.9,-6521.3,-284.02,-2606.6,-2421.9,-13608.,-1697.4,-1297.3,-5150.4,-2704.6,-5686.6,0.14307E+06,63950.,48987.,45976.,89126.,30712.,0.11009E+06,31813.,48634.,14517.,20863.,25130.,0.0000,-142.21,-148.04,-23.162,-136.33,-84.820,-558.52,-451.44,-46.323,-406.39,-48.715,-546.15
1803.000000000,8937.0,1444.4,1766.0,1852.2,2122.5,1343.4,3182.0,460.30,1860.4,353.56,753.55,853.89,0.0000,-3497.1,-6542.3,-286.80,-2605.8,-2428.9,-13607.,-1696.9,-1306.9,-5154.5,-2704.9,-5691.5,39608.,17704.,13562.,12728.,24674.,8502.6,30477.,8807.2,13464.,4018.9,5775.8,6957.3,0.0000,-39.443,-41.014,-6.4122,-37.772,-23.503,-154.62,-124.99,-12.824,-112.51,-13.487,-151.20
1804.000000000,8959.9,1443.4,1769.8,1852.4,2119.7,1326.3,3159.3,462.28,1886.4,355.85,756.25,853.83,0.0000,-3467.7,-6537.7,-285.02,-2605.1,-2407.8,-13605.,-1690.7,-1296.7,-5143.8,-2702.4,-5684.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1805.000000000,8954.8,1458.6,1765.4,1861.9,2101.2,1343.4,3182.4,463.15,1888.4,359.16,755.48,855.19,0.0000,-3458.7,-6529.0,-282.99,-2604.7,-2403.9,-13604.,-1685.9,-1291.5,-5139.5,-2701.3,-5680.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1806.000000000,8938.3,1501.3,1772.4,1888.4,2098.3,1359.7,3179.6,466.45,1899.8,362.23,757.69,855.04,0.0000,-3453.9,-6521.2,-281.40,-2604.3,-2402.2,-13604.,-1682.5,-1288.1,-5136.9,-2700.9,-5677.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1807.000000000,8926.8,1504.8,1783.6,1880.5,2096.0,1340.4,3157.4,463.80,1925.2,362.12,762.61,862.57,0.0000,-3449.6,-6515.2,-280.20,-2603.6,-2400.3,-13604.,-1680.0,-1285.4,-5135.1,-2700.4,-5675.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1808.000000000,8876.1,1499.0,1790.6,1878.9,2077.4,1321.4,3160.9,458.93,1918.4,360.09,759.16,861.45,0.0000,-3445.0,-6509.2,-279.28,-2602.7,-2398.1,-13603.,-1678.3,-1283.1,-5134.2,-2699.9,-5673.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1809.000000000,8936.6,1491.0,1802.0,1862.7,2062.7,1311.2,3174.1,454.11,1912.8,361.62,750.57,862.28,0.0000,-3440.6,-6503.3,-278.54,-2601.8,-2396.0,-13602.,-1677.0,-1281.1,-5133.0,-2699.2,-5671.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1810.000000000,8974.7,1466.5,1799.8,1843.9,2090.0,1307.7,3168.3,453.45,1915.8,360.13,755.84,865.88,0.0000,-3436.3,-6498.1,-277.93,-2601.1,-2393.8,-13601.,-1676.2,-1279.4,-5132.3,-2699.0,-5670.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1811.000000000,8972.9,1461.7,1802.8,1848.0,2111.1,1322.3,3150.7,448.42,1907.3,360.75,761.24,858.63,0.0000,-3475.1,-6516.1,-281.37,-2600.5,-2419.1,-13601.,-1676.4,-1293.8,-5143.2,-2701.2,-5677.4,5548.5,2480.1,1899.8,1783.0,3456.5,1191.1,4269.4,1233.7,1886.1,562.98,809.10,974.60,0.0000,-5.5175,-5.7394,-0.89825,-5.2871,-3.2855,-21.672,-17.513,-1.7965,-15.763,-1.8890,-21.189
1812.000000000,8984.4,1458.1,1821.4,1848.8,2120.0,1322.4,3140.7,450.01,1931.1,357.62,761.76,856.38,0.0000,-3493.1,-6536.6,-284.71,-2600.0,-2428.0,-13600.,-1682.5,-1304.6,-5147.5,-2701.8,-5681.3,50681.,22654.,17353.,16287.,31572.,10880.,38998.,11269.,17228.,5142.4,7390.5,8902.3,0.0000,-50.483,-52.455,-8.2049,-48.325,-30.044,-197.93,-159.97,-16.410,-143.99,-17.255,-193.54
1813.000000000,8977.1,1447.4,1818.5,1851.4,2137.4,1288.3,3145.6,446.47,1914.4,351.43,761.32,853.10,0.0000,-3464.4,-6532.6,-283.45,-2599.5,-2407.4,-13599.,-1680.4,-1295.0,-5137.6,-2699.6,-5674.8,0.16564,0.74040E-01,0.56717E-01,0.53231E-01,0.10319,0.35559E-01,0.12746,0.36832E-01,0.56308E-01,0.16807E-01,0.24155E-01,0.29096E-01,0.0000,-0.16497E-03,-0.17145E-03,-0.26816E-04,-0.15792E-03,-0.98008E-04,-0.64682E-03,-0.52283E-03,-0.53633E-04,-0.47059E-03,-0.56391E-04,-0.63254E-03
1814.000000000,9017.8,1453.2,1818.4,1873.3,2149.3,1300.6,3137.3,444.99,1897.0,349.04,763.84,847.33,0.0000,-3498.6,-6547.6,-285.75,-2598.8,-2430.2,-13599.,-1680.0,-1308.1,-5146.1,-2701.2,-5680.3,10220.,4567.9,3499.2,3284.1,6366.3,2193.8,7863.6,2272.4,3473.9,1036.9,1490.2,1795.1,0.0000,-10.192,-10.583,-1.6545,-9.7485,-6.0540,-39.899,-32.255,-3.3089,-29.033,-3.4792,-39.024
1815.000000000,9024.3,1442.7,1802.3,1874.3,2094.5,1279.5,3141.1,452.87,1894.4,349.90,760.69,842.22,0.0000,-3471.1,-6541.7,-284.22,-2598.0,-2410.6,-13598.,-1678.3,-1298.6,-5136.7,-2699.3,-5673.5,421.56,188.43,144.34,135.47,262.61,90.494,324.37,93.736,143.30,42.773,61.473,74.047,0.0000,-0.42027,-0.43656,-0.68246E-01,-0.40202,-0.24920,-1.6455,-1.3304,-0.13649,-1.1976,-0.14350,-1.6097
1816.000000000,9020.9,1446.7,1779.4,1868.7,2081.2,1267.1,3138.9,452.92,1894.6,349.32,758.10,836.19,0.0000,-3461.7,-6532.9,-282.49,-2597.2,-2405.9,-13596.,-1677.0,-1293.5,-5133.5,-2698.5,-5670.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1817.000000000,9095.0,1449.1,1772.3,1870.1,2083.5,1263.2,3123.2,451.39,1878.8,348.39,751.35,839.75,0.0000,-3455.0,-6523.5,-281.10,-2596.4,-2403.0,-13595.,-1676.0,-1289.9,-5131.7,-2697.8,-5668.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1818.000000000,9184.5,1442.1,1779.9,1889.5,2086.9,1278.9,3149.2,450.11,1894.6,349.06,745.63,844.98,0.0000,-3492.4,-6538.5,-283.98,-2595.6,-2428.1,-13594.,-1675.6,-1304.7,-5142.0,-2699.8,-5675.1,1384.5,618.86,474.06,444.92,862.50,297.21,1065.3,307.86,470.64,140.48,201.90,243.19,0.0000,-1.3803,-1.4336,-0.22414,-1.3201,-0.81747,-5.4023,-4.3688,-0.44829,-3.9329,-0.47126,-5.2861
1819.000000000,9199.8,1422.3,1770.9,1883.2,2092.3,1258.9,3168.4,453.58,1877.7,350.89,747.54,846.30,0.0000,-3466.1,-6533.3,-282.99,-2594.8,-2409.5,-13592.,-1675.0,-1296.2,-5133.2,-2698.1,-5668.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1820.000000000,9198.3,1425.1,1769.5,1864.9,2092.8,1259.2,3159.8,458.90,1877.2,351.67,751.53,847.93,0.0000,-3457.9,-6525.4,-281.61,-2594.0,-2405.5,-13590.,-1674.6,-1291.6,-5130.5,-2697.6,-5666.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1821.000000000,9200.5,1427.7,1781.5,1867.2,2080.1,1254.9,3164.3,456.54,1885.4,353.51,749.95,851.94,0.0000,-3452.2,-6518.0,-280.44,-2593.2,-2402.8,-13589.,-1674.2,-1288.3,-5129.3,-2697.1,-5664.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1822.000000000,9085.2,1424.9,1781.9,1877.3,2073.7,1283.4,3154.2,452.98,1902.5,353.57,746.71,855.03,0.0000,-3490.0,-6534.4,-283.47,-2592.2,-2427.6,-13588.,-1674.8,-1303.1,-5140.0,-2698.9,-5672.0,5569.5,2489.5,1907.0,1789.8,3469.5,1195.6,4285.5,1238.4,1893.2,565.11,812.16,978.29,0.0000,-5.5512,-5.7649,-0.90165,-5.3092,-3.2833,-21.725,-17.571,-1.8033,-15.820,-1.8956,-21.261
1823.000000000,9102.2,1418.8,1787.5,1891.1,2083.6,1290.4,3168.2,452.61,1907.3,351.84,745.55,857.18,0.0000,-3507.0,-6552.8,-286.52,-2591.4,-2436.3,-13587.,-1674.8,-1313.5,-5143.3,-2699.6,-5674.1,2913.4,1302.2,997.53,936.22,1814.9,625.40,2241.7,647.81,990.34,295.60,424.84,511.74,0.0000,-2.9082,-3.0172,-0.47165,-2.7790,-1.7193,-11.363,-9.1904,-0.94329,-8.2749,-0.99157,-11.121
1824.000000000,9108.6,1412.4,1792.2,1883.3,2070.3,1274.9,3170.0,454.34,1895.7,352.30,742.62,859.13,0.0000,-3477.2,-6546.6,-285.03,-2590.7,-2415.1,-13586.,-1674.4,-1302.1,-5132.9,-2697.3,-5666.7,15.028,6.7172,5.1456,4.8293,9.3618,3.2260,11.564,3.3416,5.1085,1.5248,2.1914,2.6397,0.0000,-0.14996E-01,-0.15565E-01,-0.24329E-02,-0.14332E-01,-0.88508E-02,-0.58609E-01,-0.47404E-01,-0.48658E-02,-0.42683E-01,-0.51144E-02,-0.57363E-01
1825.000000000,9141.7,1411.6,1793.1,1878.2,2083.9,1270.7,3170.1,451.35,1894.4,351.27,739.58,864.42,0.0000,-3467.4,-6536.8,-283.21,-2590.0,-2410.0,-13584.,-1674.2,-1296.2,-5129.5,-2696.3,-5664.1,760.28,339.83,260.32,244.32,473.62,163.21,585.01,169.05,258.44,77.142,110.87,133.55,0.0000,-0.75822,-0.78728,-0.12308,-0.72486,-0.44713,-2.9649,-2.3980,-0.24617,-2.1593,-0.25872,-2.9019
1826.000000000,9260.8,1405.3,1785.8,1880.5,2105.0,1294.3,3162.0,446.27,1889.8,351.38,739.51,858.40,0.0000,-3460.7,-6527.1,-281.72,-2589.4,-2406.7,-13582.,-1673.8,-1292.1,-5128.1,-2695.7,-5662.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1827.000000000,9262.5,1400.4,1776.2,1873.5,2123.8,1265.6,3165.9,445.71,1896.7,350.10,738.12,860.25,0.0000,-3454.8,-6518.5,-280.56,-2588.8,-2404.0,-13581.,-1673.6,-1288.9,-5127.1,-2694.9,-5661.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1828.000000000,9272.3,1413.9,1792.3,1888.3,2172.5,1268.7,3169.5,449.34,1914.6,353.03,739.40,858.46,0.0000,-3492.5,-6533.7,-283.61,-2588.1,-2429.0,-13581.,-1673.6,-1303.8,-5137.8,-2696.6,-5669.0,1570.7,702.08,537.81,504.75,978.48,337.18,1208.6,349.26,533.93,159.37,229.05,275.90,0.0000,-1.5660,-1.6258,-0.25428,-1.4972,-0.92332,-6.1248,-4.9532,-0.50857,-4.4607,-0.53446,-5.9944
1829.000000000,9274.3,1388.2,1791.8,1882.5,2169.1,1254.3,3150.5,453.91,1932.6,354.12,742.40,854.57,0.0000,-3466.3,-6528.5,-282.72,-2587.3,-2410.0,-13579.,-1673.4,-1295.3,-5129.4,-2694.6,-5663.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1830.000000000,9245.0,1379.8,1777.3,1875.4,2170.2,1235.7,3156.0,457.65,1938.9,351.12,742.46,851.67,0.0000,-3457.9,-6520.4,-281.41,-2586.6,-2405.4,-13578.,-1673.2,-1290.7,-5127.0,-2693.8,-5661.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1831.000000000,9222.8,1389.4,1747.5,1869.4,2183.2,1227.0,3148.1,457.42,1932.6,353.88,738.90,852.90,0.0000,-3452.0,-6512.9,-280.30,-2585.8,-2402.4,-13577.,-1673.0,-1287.5,-5126.0,-2693.0,-5660.1,3.3715,1.5070,1.1544,1.0834,2.1003,0.72375,2.5943,0.74968,1.1461,0.34209,0.49164,0.59221,0.0000,-0.33553E-02,-0.34873E-02,-0.54582E-03,-0.32107E-02,-0.19738E-02,-0.13146E-01,-0.10630E-01,-0.10916E-02,-0.95738E-02,-0.11469E-02,-0.12865E-01
1832.000000000,9174.3,1393.7,1743.4,1879.4,2174.6,1248.7,3167.4,458.21,1920.8,354.75,737.71,853.91,0.0000,-3446.7,-6505.7,-279.42,-2585.1,-2399.7,-13575.,-1672.9,-1284.8,-5125.5,-2692.3,-5659.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1833.000000000,9155.2,1392.6,1745.0,1882.0,2165.7,1250.5,3181.0,460.51,1920.7,355.20,737.11,851.53,0.0000,-3441.9,-6498.9,-278.71,-2584.4,-2397.3,-13574.,-1672.7,-1282.5,-5125.0,-2691.5,-5658.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1834.000000000,9161.2,1390.5,1746.8,1903.5,2164.9,1254.5,3171.9,462.05,1906.6,353.46,740.30,847.45,0.0000,-3437.4,-6493.0,-278.11,-2583.7,-2395.2,-13573.,-1672.6,-1280.4,-5124.7,-2690.8,-5657.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1835.000000000,9175.8,1386.5,1746.8,1895.8,2171.2,1245.8,3163.3,458.75,1902.9,350.86,739.35,843.94,0.0000,-3432.9,-6488.3,-277.61,-2583.0,-2393.0,-13572.,-1672.5,-1278.6,-5124.2,-2690.3,-5657.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1836.000000000,9184.0,1379.3,1743.6,1900.4,2183.0,1226.7,3194.6,460.47,1890.7,349.36,739.11,842.22,0.0000,-3428.5,-6483.6,-277.16,-2582.3,-2390.9,-13570.,-1672.4,-1276.9,-5123.8,-2689.8,-5656.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1837.000000000,9190.1,1370.0,1744.3,1919.0,2167.6,1219.6,3228.8,462.94,1867.9,348.04,739.05,840.42,0.0000,-3424.5,-6479.3,-276.75,-2581.7,-2388.9,-13569.,-1672.3,-1275.3,-5123.5,-2689.2,-5656.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1838.000000000,9207.4,1353.7,1752.7,1918.1,2169.0,1209.8,3241.2,462.50,1854.8,346.74,740.33,841.77,0.0000,-3420.4,-6475.4,-276.36,-2581.0,-2386.9,-13568.,-1672.2,-1273.9,-5123.3,-2688.6,-5655.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1839.000000000,9236.6,1342.9,1774.1,1912.9,2153.8,1212.1,3243.1,462.44,1853.1,347.89,741.94,840.60,0.0000,-3416.4,-6471.8,-275.99,-2580.4,-2384.9,-13566.,-1672.1,-1272.5,-5123.0,-2688.1,-5655.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1840.000000000,9251.7,1352.4,1760.6,1910.3,2149.4,1207.4,3251.4,463.28,1842.3,344.54,739.54,840.16,0.0000,-3412.7,-6468.5,-275.64,-2579.8,-2383.1,-13565.,-1672.0,-1271.3,-5122.8,-2687.6,-5655.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1841.000000000,9247.1,1351.9,1763.9,1906.7,2159.3,1196.0,3227.5,456.71,1821.7,342.93,739.65,844.35,0.0000,-3409.0,-6465.4,-275.29,-2579.3,-2381.2,-13564.,-1671.9,-1270.1,-5122.5,-2687.1,-5654.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1842.000000000,9276.2,1370.8,1768.3,1909.9,2158.0,1210.4,3210.6,454.44,1826.1,347.72,740.12,848.96,0.0000,-3448.0,-6485.3,-278.89,-2578.8,-2406.7,-13563.,-1672.3,-1283.9,-5133.6,-2689.4,-5662.0,2709.2,1211.0,927.63,870.61,1687.7,581.58,2084.6,602.41,920.94,274.89,395.06,475.88,0.0000,-2.6810,-2.7924,-0.43859,-2.5727,-1.5764,-10.561,-8.5340,-0.87719,-7.6903,-0.92112,-10.331
1843.000000000,9135.0,1365.8,1756.5,1903.1,2163.4,1191.5,3179.4,454.65,1810.4,349.61,738.97,850.73,0.0000,-3423.4,-6484.3,-278.40,-2578.3,-2388.4,-13562.,-1672.1,-1278.1,-5125.4,-2687.8,-5656.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1844.000000000,9148.4,1378.4,1758.0,1900.4,2170.3,1184.6,3159.3,458.50,1807.2,355.35,732.20,845.33,0.0000,-3416.4,-6479.8,-277.38,-2577.9,-2384.4,-13560.,-1671.9,-1275.1,-5123.0,-2687.1,-5654.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1845.000000000,9121.3,1392.6,1777.8,1910.7,2062.0,1201.2,3151.8,459.00,1808.4,358.51,729.49,838.99,0.0000,-3454.3,-6497.8,-280.40,-2577.5,-2409.3,-13560.,-1672.2,-1288.5,-5133.6,-2689.1,-5661.9,2298.8,1027.5,787.12,738.74,1432.1,493.49,1768.9,511.16,781.45,233.25,335.22,403.80,0.0000,-2.2761,-2.3696,-0.37216,-2.1834,-1.3370,-8.9600,-7.2397,-0.74432,-6.5249,-0.78153,-8.7647
1846.000000000,8937.8,1402.2,1777.6,1907.9,2087.5,1205.9,3144.1,454.83,1804.6,355.98,725.64,837.95,0.0000,-3471.6,-6518.0,-283.43,-2577.2,-2418.0,-13559.,-1672.2,-1298.7,-5136.7,-2689.8,-5664.1,1476.5,659.97,505.55,474.48,919.79,316.96,1136.1,328.31,501.91,149.81,215.31,259.35,0.0000,-1.4643,-1.5229,-0.23903,-1.4034,-0.85982,-5.7545,-4.6495,-0.47806,-4.1908,-0.50198,-5.6291
1847.000000000,8792.9,1410.9,1782.1,1896.1,2090.2,1186.1,3168.3,452.65,1802.1,358.14,718.08,837.61,0.0000,-3443.0,-6513.6,-281.94,-2576.9,-2397.2,-13557.,-1672.0,-1289.0,-5126.3,-2687.6,-5656.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1848.000000000,8867.0,1408.8,1818.0,1890.4,2098.5,1173.3,3166.0,451.61,1813.4,356.68,718.29,840.49,0.0000,-3434.2,-6505.5,-280.12,-2576.5,-2392.4,-13556.,-1671.8,-1284.0,-5123.2,-2686.7,-5654.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1849.000000000,8893.0,1412.3,1808.7,1877.9,2103.8,1161.9,3174.3,451.27,1806.8,355.10,716.36,839.35,0.0000,-3428.5,-6497.5,-278.65,-2576.1,-2389.4,-13555.,-1671.6,-1280.6,-5121.9,-2686.0,-5653.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1850.000000000,8894.5,1406.5,1806.4,1871.7,2093.4,1156.6,3175.2,454.37,1801.3,353.37,714.62,843.28,0.0000,-3423.4,-6490.3,-277.51,-2575.6,-2386.9,-13554.,-1671.4,-1277.8,-5121.1,-2685.4,-5652.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1851.000000000,8899.6,1394.2,1810.4,1885.4,2081.6,1155.9,3195.1,457.27,1795.8,351.96,714.85,841.38,0.0000,-3418.8,-6483.8,-276.62,-2575.0,-2384.6,-13553.,-1671.3,-1275.5,-5120.5,-2684.8,-5652.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1852.000000000,8853.2,1399.6,1833.0,1898.4,2059.4,1164.7,3197.9,457.89,1803.2,346.88,715.34,835.57,0.0000,-3414.5,-6478.0,-275.92,-2574.4,-2382.4,-13553.,-1671.2,-1273.5,-5120.2,-2684.3,-5651.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1853.000000000,8733.1,1395.5,1829.8,1906.5,2062.0,1159.3,3184.0,458.91,1810.8,341.84,715.69,830.97,0.0000,-3410.4,-6472.9,-275.34,-2573.8,-2380.3,-13552.,-1671.0,-1271.7,-5120.0,-2683.6,-5651.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1854.000000000,8725.9,1389.2,1825.7,1897.3,2079.2,1169.3,3160.9,461.41,1807.3,339.67,707.69,830.54,0.0000,-3406.5,-6468.3,-274.85,-2573.3,-2378.2,-13552.,-1670.9,-1270.1,-5119.7,-2682.9,-5650.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1855.000000000,8722.0,1383.1,1791.0,1879.7,2077.8,1170.0,3183.9,463.21,1796.6,341.17,702.57,836.56,0.0000,-3402.8,-6464.0,-274.42,-2572.8,-2376.2,-13551.,-1670.8,-1268.7,-5119.3,-2682.2,-5650.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1856.000000000,8725.9,1383.1,1778.8,1845.4,2068.2,1181.8,3200.9,462.52,1807.4,341.32,700.07,834.62,0.0000,-3399.2,-6459.9,-274.03,-2572.3,-2374.3,-13550.,-1670.8,-1267.3,-5118.9,-2681.6,-5650.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1857.000000000,8620.3,1384.3,1780.3,1836.3,2061.2,1200.3,3202.9,459.63,1807.8,342.27,704.93,832.69,0.0000,-3395.8,-6456.2,-273.67,-2571.7,-2372.4,-13549.,-1670.7,-1266.0,-5118.5,-2681.1,-5649.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1858.000000000,8631.6,1375.5,1776.4,1827.8,2059.1,1179.3,3197.5,460.05,1819.0,344.31,704.51,832.43,0.0000,-3392.6,-6453.0,-273.33,-2571.2,-2370.6,-13549.,-1670.6,-1264.8,-5118.2,-2680.6,-5649.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1859.000000000,8572.7,1373.4,1783.1,1831.7,2183.2,1176.8,3185.6,459.73,1825.0,341.80,704.10,832.01,0.0000,-3389.4,-6450.0,-273.02,-2570.6,-2368.8,-13548.,-1670.5,-1263.9,-5117.9,-2680.1,-5649.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1860.000000000,8532.1,1378.1,1786.9,1835.9,2290.2,1197.1,3170.1,463.87,1837.4,338.85,701.33,823.32,0.0000,-3428.6,-6470.2,-276.65,-2570.1,-2394.3,-13547.,-1670.9,-1277.3,-5129.1,-2682.1,-5656.7,3041.2,1359.3,1041.3,977.29,1894.5,652.84,2340.1,676.23,1033.8,308.57,443.47,534.19,0.0000,-2.9975,-3.1247,-0.49234,-2.8806,-1.7540,-11.843,-9.5666,-0.98468,-8.6301,-1.0331,-11.586
1861.000000000,8543.8,1380.6,1786.3,1833.5,2283.0,1183.0,3141.4,459.67,1808.6,336.65,706.18,826.59,0.0000,-3404.5,-6469.4,-276.22,-2569.6,-2376.0,-13546.,-1670.7,-1272.3,-5121.0,-2680.3,-5651.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1862.000000000,8556.8,1372.2,1767.1,1842.7,2301.2,1183.1,3152.9,458.56,1799.9,336.87,699.79,828.78,0.0000,-3397.9,-6465.0,-275.24,-2569.2,-2372.1,-13545.,-1670.5,-1269.6,-5118.7,-2679.4,-5649.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1863.000000000,8600.6,1365.5,1755.9,1837.6,2129.9,1180.6,3143.5,457.38,1793.7,338.38,698.80,823.47,0.0000,-3393.5,-6460.2,-274.36,-2568.9,-2369.7,-13544.,-1670.4,-1267.4,-5117.5,-2678.7,-5648.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1864.000000000,8588.3,1373.3,1759.9,1846.2,2110.6,1195.6,3147.5,458.95,1786.7,341.18,695.02,821.99,0.0000,-3432.0,-6478.7,-277.59,-2568.6,-2395.1,-13543.,-1670.5,-1280.4,-5128.3,-2680.6,-5656.0,1368.1,611.53,468.45,439.65,852.29,293.69,1052.7,304.21,465.07,138.82,199.51,240.31,0.0000,-1.3487,-1.4053,-0.22149,-1.2958,-0.78819,-5.3260,-4.3024,-0.44298,-3.8822,-0.46467,-5.2111
1865.000000000,8515.7,1367.3,1753.3,1833.8,2108.9,1192.6,3156.4,456.91,1773.9,341.78,692.82,826.92,0.0000,-3407.3,-6476.2,-276.86,-2568.1,-2376.6,-13541.,-1670.3,-1274.3,-5120.0,-2678.8,-5650.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1866.000000000,8400.3,1347.6,1786.3,1837.3,2110.0,1190.9,3165.8,459.06,1770.3,342.77,697.00,834.07,0.0000,-3400.2,-6470.4,-275.70,-2567.6,-2372.7,-13540.,-1670.2,-1271.0,-5117.6,-2677.9,-5648.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1867.000000000,8413.3,1338.1,1802.1,1835.7,2114.6,1185.4,3150.5,454.51,1762.4,339.97,701.02,836.36,0.0000,-3395.3,-6464.4,-274.69,-2567.1,-2370.2,-13538.,-1670.0,-1268.6,-5116.5,-2677.2,-5647.6,2.6120,1.1675,0.89434,0.83937,1.6272,0.56071,2.0098,0.58079,0.88789,0.26503,0.38089,0.45880,0.0000,-0.25715E-02,-0.26814E-02,-0.42286E-03,-0.24722E-02,-0.15001E-02,-0.10166E-01,-0.82122E-02,-0.84571E-03,-0.74115E-02,-0.88691E-03,-0.99473E-02
1868.000000000,8248.3,1339.5,1783.3,1829.3,2121.9,1165.1,3149.0,454.55,1749.4,342.70,700.01,833.40,0.0000,-3391.0,-6458.6,-273.88,-2566.5,-2368.0,-13537.,-1669.9,-1266.7,-5115.8,-2676.7,-5647.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1869.000000000,8095.0,1348.4,1760.9,1839.5,2116.1,1159.7,3138.4,454.62,1748.3,341.69,703.65,829.69,0.0000,-3386.9,-6453.3,-273.24,-2566.0,-2366.0,-13536.,-1669.8,-1265.0,-5115.3,-2676.1,-5646.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1870.000000000,8060.9,1358.3,1765.5,1840.4,2112.1,1176.7,3139.5,453.14,1768.8,341.51,705.11,825.69,0.0000,-3425.4,-6471.5,-276.64,-2565.5,-2391.4,-13535.,-1671.0,-1277.9,-5126.4,-2678.1,-5654.2,9693.6,4332.8,3319.1,3115.1,6038.7,2080.9,7458.9,2155.4,3295.1,983.56,1413.5,1702.7,0.0000,-9.5452,-9.9474,-1.5693,-9.1746,-5.5710,-37.720,-30.471,-3.1386,-27.505,-3.2911,-36.911
1871.000000000,8063.7,1355.2,1769.0,1839.3,2116.9,1175.8,3117.4,449.21,1771.0,342.82,704.24,827.01,0.0000,-3443.2,-6492.3,-279.99,-2565.1,-2400.2,-13535.,-1671.1,-1288.2,-5129.7,-2678.7,-5656.9,3318.5,1483.3,1136.3,1066.4,2067.3,712.37,2553.5,737.89,1128.1,336.71,483.92,582.90,0.0000,-3.2733,-3.4074,-0.53724,-3.1431,-1.9099,-12.913,-10.431,-1.0745,-9.4159,-1.1267,-12.636
1872.000000000,8146.8,1336.8,1753.5,1832.0,2109.1,1163.4,3117.5,449.72,1779.2,342.28,700.03,829.30,0.0000,-3414.9,-6488.5,-278.73,-2564.7,-2379.6,-13533.,-1670.7,-1279.4,-5119.5,-2676.4,-5650.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1873.000000000,8160.9,1324.8,1758.4,1827.9,2095.6,1156.0,3110.7,455.29,1772.1,343.34,701.45,829.47,0.0000,-3406.3,-6480.8,-277.08,-2564.1,-2374.7,-13532.,-1670.3,-1274.8,-5116.4,-2675.3,-5647.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1874.000000000,8167.9,1324.3,1757.5,1823.8,2183.9,1142.9,3112.3,456.32,1767.3,341.41,694.26,831.68,0.0000,-3400.5,-6473.0,-275.71,-2563.5,-2371.7,-13530.,-1669.9,-1271.8,-5115.0,-2674.4,-5646.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1875.000000000,8168.4,1323.3,1751.6,1818.2,2307.5,1141.6,3112.1,455.91,1780.2,343.73,691.64,823.06,0.0000,-3395.4,-6466.0,-274.64,-2563.0,-2369.2,-13529.,-1669.7,-1269.6,-5114.1,-2673.6,-5645.6,40.942,18.300,14.018,13.157,25.505,8.7889,31.504,9.1037,13.917,4.1542,5.9703,7.1915,0.0000,-0.40311E-01,-0.42009E-01,-0.66281E-02,-0.38742E-01,-0.23452E-01,-0.15929,-0.12865,-0.13256E-01,-0.11616,-0.13896E-01,-0.15586
1876.000000000,8364.3,1323.3,1755.2,1827.1,2312.6,1159.3,3124.2,455.03,1774.5,344.66,693.75,824.69,0.0000,-3433.3,-6482.9,-277.75,-2562.5,-2394.2,-13528.,-1671.5,-1283.1,-5125.3,-2675.3,-5653.3,14321.,6401.1,4903.4,4602.0,8921.2,3074.2,11019.,3184.3,4868.0,1453.0,2088.3,2515.4,0.0000,-14.119,-14.698,-2.3184,-13.559,-8.2197,-55.715,-44.997,-4.6368,-40.631,-4.8605,-54.515
1877.000000000,8393.3,1323.3,1754.0,1829.7,2311.4,1162.9,3130.9,456.08,1764.6,342.82,690.62,825.26,0.0000,-3450.5,-6502.3,-280.87,-2562.2,-2402.7,-13528.,-1676.4,-1293.2,-5129.6,-2675.7,-5657.2,41223.,18426.,14115.,13247.,25680.,8849.2,31720.,9166.2,14013.,4182.7,6011.2,7240.9,0.0000,-40.711,-42.334,-6.6736,-39.056,-23.693,-160.38,-129.53,-13.347,-116.96,-13.991,-156.92
1878.000000000,8430.5,1321.4,1752.4,1835.3,2315.2,1164.5,3126.8,455.50,1748.0,341.04,689.24,822.69,0.0000,-3464.5,-6520.4,-283.39,-2562.0,-2409.2,-13527.,-1696.6,-1301.5,-5135.7,-2675.8,-5664.6,0.16557E+06,74009.,56693.,53208.,0.10315E+06,35543.,0.12740E+06,36817.,56284.,16800.,24145.,29083.,0.0000,-163.81,-170.16,-26.805,-156.99,-95.263,-644.15,-520.33,-53.610,-469.78,-56.198,-630.29
1879.000000000,8443.2,1315.8,1761.7,1847.3,2316.5,1163.2,3145.1,458.89,1754.6,341.59,687.20,828.80,0.0000,-3477.4,-6536.7,-285.38,-2561.8,-2415.1,-13527.,-1691.1,-1308.7,-5138.5,-2675.8,-5668.1,12041.,5382.3,4122.9,3869.5,7501.2,2584.9,9265.4,2677.5,4093.2,1221.8,1755.9,2115.1,0.0000,-11.935,-12.386,-1.9494,-11.426,-6.9342,-46.851,-37.845,-3.8988,-34.165,-4.0869,-45.841
1880.000000000,8456.9,1307.6,1751.4,1850.6,2326.4,1168.0,3168.0,462.22,1741.1,344.66,688.24,835.32,0.0000,-3446.5,-6528.1,-283.04,-2562.0,-2394.3,-13526.,-1685.1,-1295.7,-5127.0,-2673.4,-5660.2,567.90,253.84,194.45,182.50,353.78,121.91,436.98,126.28,193.05,57.622,82.813,99.753,0.0000,-0.56304,-0.58441,-0.91938E-01,-0.53905,-0.32693,-2.2106,-1.7852,-0.18388,-1.6114,-0.19274,-2.1626
1881.000000000,8377.1,1342.4,1761.1,1837.5,2329.9,1185.8,3164.5,461.51,1739.5,340.46,694.10,834.39,0.0000,-3480.9,-6540.3,-284.60,-2562.3,-2417.8,-13527.,-1680.9,-1307.6,-5134.0,-2675.2,-5664.1,3573.4,1597.2,1223.5,1148.3,2226.1,767.09,2749.6,794.57,1214.7,362.58,521.08,627.67,0.0000,-3.5508,-3.6802,-0.57850,-3.3958,-2.0650,-13.916,-11.235,-1.1570,-10.140,-1.2133,-13.610
1882.000000000,8311.1,1311.9,1768.5,1823.6,2310.1,1164.5,3126.9,456.31,1718.9,340.35,703.03,840.61,0.0000,-3453.0,-6532.6,-282.55,-2562.2,-2398.0,-13527.,-1677.4,-1296.1,-5123.7,-2673.2,-5656.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1883.000000000,8451.2,1311.7,1772.8,1824.1,2306.4,1152.3,3095.8,453.87,1714.3,340.62,696.73,841.34,0.0000,-3443.3,-6521.8,-280.44,-2561.8,-2392.6,-13526.,-1674.9,-1289.7,-5120.1,-2672.2,-5652.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1884.000000000,8509.0,1302.9,1768.2,1825.1,2316.9,1146.5,3093.6,452.50,1714.8,342.02,695.31,845.11,0.0000,-3435.6,-6510.8,-278.76,-2561.3,-2388.8,-13525.,-1673.1,-1285.1,-5117.9,-2671.2,-5649.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1885.000000000,8506.2,1323.1,1765.6,1818.9,2331.3,1139.1,3090.5,449.92,1705.5,340.17,698.92,848.44,0.0000,-3429.4,-6500.8,-277.46,-2561.1,-2385.6,-13524.,-1671.9,-1281.3,-5116.3,-2671.0,-5647.6,10.334,4.6193,3.5385,3.3210,6.4379,2.2185,7.9520,2.2979,3.5130,1.0486,1.5070,1.8153,0.0000,-0.10240E-01,-0.10633E-01,-0.16731E-02,-0.98064E-02,-0.59473E-02,-0.40244E-01,-0.32498E-01,-0.33461E-02,-0.29327E-01,-0.35072E-02,-0.39369E-01
1886.000000000,8617.3,1329.8,1780.6,1828.5,2343.5,1146.9,3075.3,448.78,1719.4,339.84,697.05,848.10,0.0000,-3466.7,-6515.3,-280.41,-2560.9,-2410.1,-13524.,-1672.2,-1295.4,-5126.6,-2672.9,-5654.5,8593.0,3840.9,2942.2,2761.4,5353.1,1844.6,6612.0,1910.7,2921.0,871.89,1253.1,1509.4,0.0000,-8.5249,-8.8433,-1.3911,-8.1576,-4.9544,-33.460,-27.022,-2.7823,-24.385,-2.9163,-32.735
1887.000000000,8631.5,1338.9,1778.2,1822.4,2344.9,1146.9,3080.7,448.72,1726.0,339.62,694.83,845.63,0.0000,-3440.0,-6509.7,-279.45,-2560.5,-2390.8,-13523.,-1671.3,-1286.7,-5117.8,-2670.8,-5648.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1888.000000000,8666.1,1332.3,1774.7,1821.1,2347.0,1155.2,3086.4,452.49,1716.4,338.68,698.64,848.36,0.0000,-3431.2,-6501.1,-278.09,-2559.9,-2386.0,-13522.,-1670.6,-1281.8,-5115.0,-2670.0,-5646.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1889.000000000,8737.8,1331.0,1775.9,1826.0,2351.7,1159.4,3085.3,449.41,1721.7,335.92,700.40,849.45,0.0000,-3424.9,-6493.0,-276.94,-2559.3,-2382.8,-13521.,-1670.0,-1278.2,-5113.5,-2669.4,-5644.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1890.000000000,8742.9,1338.5,1775.6,1832.3,2366.5,1162.4,3085.7,442.78,1714.6,333.25,697.75,846.47,0.0000,-3419.2,-6485.7,-276.03,-2558.7,-2379.9,-13520.,-1669.6,-1275.3,-5112.6,-2668.9,-5643.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1891.000000000,8813.8,1332.7,1769.3,1829.3,2366.4,1155.0,3082.9,444.55,1707.4,332.64,698.31,844.52,0.0000,-3413.9,-6478.5,-275.30,-2558.1,-2377.2,-13519.,-1669.3,-1272.8,-5111.8,-2668.5,-5643.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1892.000000000,8847.7,1333.7,1745.9,1829.9,2346.0,1148.0,3074.5,450.76,1709.1,333.04,690.27,843.99,0.0000,-3409.0,-6472.0,-274.70,-2557.5,-2374.6,-13518.,-1669.0,-1270.6,-5111.2,-2668.1,-5642.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1893.000000000,8692.8,1337.6,1742.7,1842.0,2350.9,1138.1,3067.0,448.93,1700.5,333.20,687.39,846.66,0.0000,-3404.4,-6466.2,-274.18,-2556.9,-2372.1,-13517.,-1668.8,-1268.8,-5110.5,-2667.7,-5641.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1894.000000000,8705.4,1333.5,1744.9,1813.3,2351.9,1141.3,3061.9,448.32,1700.4,332.70,685.08,844.13,0.0000,-3400.0,-6461.2,-273.73,-2556.3,-2369.7,-13516.,-1668.7,-1267.2,-5109.9,-2667.6,-5641.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1895.000000000,8693.0,1316.7,1762.7,1809.4,2343.2,1144.1,3042.1,444.87,1692.3,331.56,685.39,843.00,0.0000,-3395.8,-6456.7,-273.32,-2555.7,-2367.4,-13515.,-1668.5,-1265.7,-5109.3,-2667.4,-5640.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1896.000000000,8700.0,1304.7,1769.9,1816.2,2343.3,1156.7,3035.5,443.73,1676.0,328.45,684.11,838.37,0.0000,-3391.9,-6452.4,-272.95,-2555.2,-2365.2,-13514.,-1668.4,-1264.3,-5108.7,-2667.1,-5640.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1897.000000000,8698.7,1314.6,1764.9,1836.3,2347.7,1170.2,3035.2,442.88,1693.0,324.63,680.27,840.14,0.0000,-3388.3,-6448.3,-272.59,-2554.6,-2363.0,-13514.,-1668.3,-1263.0,-5108.0,-2666.6,-5639.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1898.000000000,8709.3,1319.4,1751.3,1834.8,2289.2,1161.3,3011.0,442.18,1703.8,324.06,682.88,835.01,0.0000,-3384.8,-6444.4,-272.25,-2554.1,-2360.8,-13513.,-1668.2,-1261.7,-5107.4,-2666.1,-5638.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1899.000000000,8719.1,1322.9,1744.2,1842.1,2201.9,1153.2,3009.3,440.87,1693.0,322.30,679.46,831.61,0.0000,-3381.3,-6440.9,-271.92,-2553.6,-2358.7,-13512.,-1668.1,-1260.4,-5106.8,-2665.6,-5638.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1900.000000000,8823.3,1326.9,1801.1,1815.2,2182.7,1153.6,3007.3,435.55,1695.1,318.17,680.92,828.89,0.0000,-3377.8,-6437.5,-271.59,-2553.0,-2356.6,-13511.,-1668.0,-1259.2,-5106.2,-2665.0,-5638.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1901.000000000,8899.6,1320.5,1851.4,1804.5,2189.7,1154.7,3038.9,434.31,1691.3,317.47,680.60,826.26,0.0000,-3374.6,-6434.2,-271.27,-2552.5,-2354.5,-13510.,-1667.9,-1258.1,-5105.6,-2664.4,-5637.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1902.000000000,9084.0,1319.1,1838.3,1799.5,2176.5,1138.4,3047.2,434.43,1683.2,314.29,680.73,824.07,0.0000,-3371.3,-6431.1,-270.96,-2552.0,-2352.5,-13509.,-1667.8,-1257.0,-5105.1,-2663.8,-5637.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1903.000000000,9086.7,1311.5,1825.6,1786.6,2166.0,1121.4,3032.8,433.29,1672.0,311.66,686.01,829.53,0.0000,-3368.0,-6428.2,-270.65,-2551.5,-2350.6,-13509.,-1667.7,-1256.0,-5104.6,-2663.3,-5637.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1904.000000000,9055.8,1298.6,1823.7,1778.6,2158.3,1113.2,3028.5,435.71,1678.7,309.34,691.31,826.33,0.0000,-3364.8,-6425.4,-270.35,-2551.0,-2348.7,-13508.,-1667.6,-1255.1,-5104.1,-2662.7,-5636.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1905.000000000,8956.1,1290.5,1826.4,1770.5,2162.4,1108.6,3025.0,434.43,1674.7,308.31,693.36,816.18,0.0000,-3361.7,-6422.6,-270.03,-2550.5,-2346.9,-13507.,-1667.6,-1254.2,-5103.7,-2662.2,-5636.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1906.000000000,8700.1,1304.1,1818.6,1760.4,2168.2,1109.3,3031.2,431.53,1683.7,306.72,688.44,813.39,0.0000,-3358.7,-6420.0,-269.70,-2549.9,-2345.2,-13507.,-1667.5,-1253.4,-5103.3,-2661.5,-5636.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1907.000000000,8658.3,1297.9,1820.5,1760.4,2178.3,1108.5,3007.7,430.95,1685.3,305.00,682.48,810.23,0.0000,-3355.9,-6417.6,-269.38,-2549.4,-2343.5,-13506.,-1667.4,-1252.6,-5102.8,-2660.9,-5636.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1908.000000000,8555.9,1300.6,1824.1,1755.8,2174.3,1112.8,2998.3,432.72,1675.8,304.62,679.55,810.25,0.0000,-3353.0,-6415.2,-269.07,-2548.8,-2341.8,-13506.,-1667.3,-1251.9,-5102.3,-2660.3,-5635.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1909.000000000,8521.8,1292.2,1832.7,1752.9,2174.1,1096.0,3004.4,431.24,1666.4,305.16,678.81,811.32,0.0000,-3350.4,-6413.2,-268.76,-2548.3,-2340.1,-13505.,-1667.2,-1251.2,-5101.8,-2659.7,-5635.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1910.000000000,8493.4,1291.4,1831.5,1756.7,2184.7,1085.8,2976.6,433.33,1658.8,302.81,676.21,805.34,0.0000,-3347.8,-6411.0,-268.45,-2547.7,-2338.5,-13504.,-1667.2,-1250.5,-5101.4,-2659.2,-5635.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1911.000000000,8487.1,1299.8,1819.2,1740.3,2184.2,1077.6,2946.1,437.21,1662.3,301.97,671.74,800.38,0.0000,-3345.2,-6408.8,-268.15,-2547.1,-2336.8,-13503.,-1667.1,-1249.9,-5101.0,-2658.6,-5634.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1912.000000000,8477.7,1300.9,1838.2,1730.8,2167.2,1078.4,2937.0,437.98,1669.7,300.41,668.90,795.21,0.0000,-3342.7,-6406.6,-267.86,-2546.6,-2335.1,-13502.,-1667.0,-1249.3,-5100.6,-2658.1,-5634.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1913.000000000,8469.8,1305.6,1848.1,1742.2,2154.0,1107.3,2935.4,436.50,1673.3,300.64,667.66,794.27,0.0000,-3382.0,-6427.4,-271.49,-2546.2,-2360.7,-13502.,-1668.1,-1260.0,-5111.8,-2660.0,-5642.4,8141.5,3639.1,2787.6,2616.3,5071.8,1747.7,6264.6,1810.3,2767.5,826.08,1187.2,1430.1,0.0000,-7.9527,-8.3044,-1.3180,-7.6753,-4.6076,-31.640,-25.556,-2.6361,-23.097,-2.7600,-30.980
1914.000000000,8474.1,1299.8,1849.5,1713.6,2157.5,1109.8,2914.4,434.48,1655.3,303.39,662.52,795.66,0.0000,-3358.5,-6427.3,-271.05,-2545.7,-2342.5,-13500.,-1667.7,-1256.2,-5103.7,-2658.0,-5637.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1915.000000000,8468.4,1302.4,1838.6,1722.3,2156.1,1123.0,2900.5,432.53,1655.4,304.44,663.64,797.13,0.0000,-3352.4,-6423.5,-270.08,-2545.3,-2338.7,-13499.,-1667.4,-1254.0,-5101.2,-2657.0,-5635.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1916.000000000,8502.1,1306.2,1832.1,1742.3,2139.9,1114.2,2894.6,432.03,1646.2,307.72,664.29,791.64,0.0000,-3348.5,-6419.2,-269.21,-2544.9,-2336.4,-13497.,-1667.2,-1252.5,-5100.1,-2656.3,-5634.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1917.000000000,8593.6,1307.3,1826.7,1756.1,2136.9,1116.8,2903.6,438.25,1657.7,307.39,669.24,790.58,0.0000,-3345.1,-6415.3,-268.51,-2544.5,-2334.5,-13496.,-1667.0,-1251.3,-5099.4,-2655.8,-5633.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1918.000000000,8599.3,1300.1,1822.2,1759.2,2130.1,1122.8,2904.0,438.84,1664.9,308.52,667.73,792.08,0.0000,-3341.9,-6411.7,-267.94,-2544.0,-2332.7,-13494.,-1666.8,-1250.2,-5098.9,-2655.3,-5633.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1919.000000000,8622.0,1295.2,1818.1,1746.9,2123.5,1127.2,2924.8,433.53,1654.4,307.95,666.24,790.00,0.0000,-3338.8,-6408.8,-267.46,-2543.6,-2331.1,-13493.,-1666.6,-1249.2,-5098.4,-2654.9,-5633.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1920.000000000,8631.4,1295.7,1819.0,1751.1,2142.4,1119.1,2920.6,430.29,1650.9,308.96,668.76,794.13,0.0000,-3335.9,-6406.4,-267.04,-2543.1,-2329.6,-13492.,-1666.5,-1248.3,-5098.0,-2654.5,-5632.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1921.000000000,8640.5,1291.1,1829.8,1745.6,2146.3,1116.6,2905.9,429.31,1644.6,308.86,671.73,797.35,0.0000,-3333.1,-6404.3,-266.66,-2542.6,-2328.1,-13490.,-1666.4,-1247.5,-5097.3,-2654.0,-5632.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1922.000000000,8642.2,1281.0,1830.2,1738.3,2136.9,1109.8,2915.4,424.86,1635.6,308.42,677.17,794.24,0.0000,-3330.3,-6402.3,-266.32,-2542.1,-2326.5,-13489.,-1666.3,-1246.8,-5096.8,-2653.5,-5632.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1923.000000000,8638.7,1298.4,1839.2,1725.7,2124.7,1109.4,2906.3,429.78,1635.1,308.59,675.33,788.76,0.0000,-3327.6,-6400.3,-266.00,-2541.6,-2325.1,-13488.,-1666.2,-1246.2,-5096.3,-2653.0,-5631.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1924.000000000,8638.5,1302.2,1835.8,1723.2,2106.3,1103.3,2904.6,432.01,1626.9,306.44,677.39,787.39,0.0000,-3325.0,-6398.1,-265.70,-2541.1,-2323.6,-13487.,-1666.1,-1245.5,-5095.9,-2652.4,-5631.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1925.000000000,8637.3,1312.0,1826.8,1713.4,2105.6,1095.6,2896.2,432.05,1619.6,304.68,681.75,784.00,0.0000,-3322.5,-6396.0,-265.42,-2540.6,-2322.1,-13486.,-1666.1,-1244.9,-5095.4,-2651.8,-5631.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1926.000000000,8621.7,1310.2,1827.2,1698.6,2106.3,1087.0,2898.7,435.87,1626.3,301.85,679.84,778.95,0.0000,-3320.1,-6393.9,-265.16,-2540.1,-2320.7,-13485.,-1666.0,-1244.2,-5095.1,-2651.3,-5630.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1927.000000000,8598.0,1292.9,1818.5,1711.4,2103.1,1085.1,2903.7,439.61,1622.6,301.92,677.57,771.16,0.0000,-3317.7,-6391.9,-264.91,-2539.6,-2319.2,-13483.,-1665.9,-1243.6,-5095.0,-2650.8,-5630.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1928.000000000,8454.6,1291.1,1805.5,1704.5,2104.2,1088.0,2911.1,441.79,1602.6,300.90,675.02,766.93,0.0000,-3315.3,-6390.1,-264.67,-2539.1,-2317.8,-13482.,-1665.8,-1243.0,-5094.9,-2650.3,-5629.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1929.000000000,8384.1,1289.9,1813.1,1694.7,2122.7,1085.3,2920.1,441.47,1589.1,296.36,674.70,764.29,0.0000,-3312.9,-6388.3,-264.44,-2538.8,-2316.3,-13481.,-1665.8,-1242.4,-5094.8,-2649.8,-5629.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1930.000000000,8450.7,1281.7,1804.1,1696.4,2126.4,1094.0,2900.2,437.64,1595.2,294.70,672.89,760.72,0.0000,-3352.1,-6409.3,-268.12,-2538.6,-2342.1,-13481.,-1666.3,-1251.8,-5106.0,-2651.8,-5636.8,4400.4,1966.9,1506.7,1414.1,2741.2,944.62,3386.0,978.46,1495.8,446.49,641.68,772.93,0.0000,-4.2716,-4.4694,-0.71238,-4.1370,-2.4724,-17.078,-13.796,-1.4248,-12.481,-1.4909,-16.732
1931.000000000,8508.0,1276.9,1797.3,1705.7,2125.4,1078.1,2890.5,436.57,1581.4,294.83,669.07,754.86,0.0000,-3328.8,-6409.3,-267.76,-2538.5,-2324.2,-13479.,-1666.1,-1248.5,-5097.8,-2650.0,-5631.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1932.000000000,8515.7,1262.6,1808.7,1708.5,2126.1,1067.0,2890.1,434.47,1580.0,294.06,667.25,754.91,0.0000,-3322.9,-6405.8,-266.85,-2538.3,-2320.5,-13478.,-1665.9,-1246.7,-5095.4,-2649.1,-5629.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1933.000000000,8487.3,1267.8,1818.0,1686.0,2127.4,1061.7,2893.2,438.42,1604.0,298.29,667.79,752.92,0.0000,-3319.3,-6401.8,-266.04,-2538.1,-2318.3,-13477.,-1665.7,-1245.5,-5094.3,-2648.4,-5628.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1934.000000000,8410.3,1270.7,1813.2,1665.2,2123.5,1057.2,2900.2,438.30,1612.0,298.76,669.52,749.02,0.0000,-3316.3,-6398.2,-265.39,-2537.8,-2316.5,-13476.,-1665.6,-1244.4,-5093.4,-2647.7,-5628.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1935.000000000,8413.4,1271.5,1798.6,1663.1,2123.1,1049.9,2885.9,435.21,1616.7,295.46,670.60,752.47,0.0000,-3313.4,-6395.1,-264.88,-2537.3,-2314.8,-13475.,-1665.5,-1243.5,-5092.6,-2647.2,-5627.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1936.000000000,8462.8,1284.8,1791.2,1669.4,2120.2,1042.0,2882.1,434.32,1613.2,294.12,667.29,748.89,0.0000,-3310.8,-6392.1,-264.46,-2536.8,-2313.2,-13474.,-1665.3,-1242.7,-5092.1,-2646.6,-5627.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1937.000000000,8665.5,1277.6,1782.6,1683.0,2102.0,1033.8,2891.9,434.50,1603.4,292.66,665.53,749.09,0.0000,-3308.2,-6389.4,-264.10,-2536.2,-2311.6,-13473.,-1665.3,-1241.9,-5091.6,-2646.1,-5626.8,671.18,300.01,229.81,215.69,418.12,144.08,516.45,149.24,228.16,68.102,97.874,117.89,0.0000,-0.64989,-0.68071,-0.10866,-0.63018,-0.37519,-2.6032,-2.1032,-0.21732,-1.9035,-0.22735,-2.5514
1938.000000000,8654.5,1282.5,1784.0,1699.7,2085.3,1047.7,2875.6,438.18,1593.9,293.46,665.87,749.34,0.0000,-3347.2,-6409.7,-267.69,-2535.7,-2337.3,-13473.,-1665.6,-1251.4,-5102.6,-2648.0,-5634.3,2656.7,1187.5,909.64,853.73,1655.0,570.30,2044.2,590.73,903.09,269.56,387.41,466.65,0.0000,-2.5758,-2.6954,-0.43009,-2.4960,-1.4886,-10.303,-8.3242,-0.86018,-7.5345,-0.89991,-10.098
1939.000000000,8648.9,1294.1,1778.3,1699.8,2076.2,1040.4,2879.0,440.39,1575.5,291.76,668.27,750.59,0.0000,-3323.9,-6409.2,-267.26,-2535.4,-2319.3,-13472.,-1665.4,-1248.0,-5094.3,-2646.1,-5628.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1940.000000000,8591.7,1295.0,1777.8,1684.1,2075.6,1030.4,2875.3,438.04,1565.4,291.92,666.78,753.88,0.0000,-3318.0,-6405.2,-266.31,-2535.1,-2315.7,-13470.,-1665.3,-1246.0,-5091.8,-2645.2,-5627.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1941.000000000,8565.8,1278.4,1764.4,1689.7,2077.3,1032.5,2876.8,435.59,1574.5,290.82,665.68,753.21,0.0000,-3314.3,-6400.9,-265.47,-2534.6,-2313.6,-13470.,-1665.1,-1244.6,-5090.8,-2644.5,-5626.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1942.000000000,8561.4,1269.1,1743.1,1684.6,1974.5,1060.4,2874.4,434.32,1597.2,290.50,660.27,751.70,0.0000,-3352.6,-6419.7,-268.72,-2534.2,-2339.0,-13469.,-1668.6,-1254.6,-5102.2,-2646.4,-5634.3,27214.,12164.,9318.0,8745.2,16953.,5841.9,20940.,6051.2,9250.8,2761.3,3968.4,4780.1,0.0000,-26.404,-27.612,-4.4057,-25.574,-15.240,-105.50,-85.249,-8.8113,-77.176,-9.2173,-103.43
1943.000000000,8624.3,1275.2,1715.8,1669.9,2014.2,1051.5,2883.2,431.63,1593.7,291.69,657.71,751.87,0.0000,-3328.7,-6417.9,-268.05,-2533.8,-2320.8,-13468.,-1667.6,-1250.4,-5094.2,-2644.5,-5629.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1944.000000000,8607.9,1271.6,1726.0,1658.1,1996.7,1043.4,2869.6,430.22,1591.9,290.54,657.71,753.54,0.0000,-3322.3,-6413.0,-266.93,-2533.4,-2317.0,-13467.,-1666.8,-1248.0,-5091.6,-2643.6,-5627.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1945.000000000,8795.8,1269.8,1715.9,1655.6,1992.1,1038.3,2865.1,428.58,1593.4,289.25,656.16,754.33,0.0000,-3318.2,-6408.0,-265.98,-2532.9,-2314.7,-13466.,-1666.1,-1246.3,-5090.3,-2642.8,-5626.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1946.000000000,8841.0,1283.5,1721.3,1653.5,1981.9,1033.2,2882.0,428.51,1587.6,289.49,654.22,751.43,0.0000,-3314.6,-6403.3,-265.24,-2532.4,-2312.8,-13465.,-1665.6,-1244.9,-5089.4,-2642.2,-5625.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1947.000000000,8846.0,1288.3,1717.1,1647.8,1983.9,1034.7,2873.3,427.79,1586.6,288.81,650.14,750.16,0.0000,-3311.3,-6399.1,-264.67,-2531.9,-2311.0,-13464.,-1665.2,-1243.7,-5088.6,-2641.6,-5624.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1948.000000000,8994.0,1289.5,1711.0,1646.2,1981.9,1032.8,2865.6,427.87,1577.6,288.01,650.14,749.84,0.0000,-3308.2,-6395.4,-264.25,-2531.4,-2309.3,-13463.,-1664.9,-1242.6,-5087.9,-2641.0,-5623.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1949.000000000,9060.6,1294.3,1716.1,1638.2,1982.4,1051.5,2877.1,427.18,1585.6,288.10,652.83,749.64,0.0000,-3346.8,-6414.9,-267.82,-2530.9,-2334.9,-13463.,-1665.9,-1252.4,-5098.9,-2643.0,-5631.5,8371.7,3742.0,2866.4,2690.3,5215.2,1797.1,6441.7,1861.5,2845.8,849.43,1220.8,1470.5,0.0000,-8.1149,-8.4866,-1.3553,-7.8632,-4.6770,-32.433,-26.213,-2.7106,-23.739,-2.8348,-31.810
1950.000000000,8956.9,1296.0,1713.7,1641.0,1989.5,1068.6,2880.1,425.07,1599.1,287.78,650.21,748.44,0.0000,-3364.7,-6436.3,-271.31,-2530.7,-2344.1,-13462.,-1690.7,-1261.3,-5107.3,-2643.6,-5640.7,0.18990E+06,84881.,65021.,61024.,0.11830E+06,40765.,0.14612E+06,42225.,64552.,19268.,27692.,33356.,0.0000,-184.40,-192.63,-30.743,-178.51,-106.26,-735.64,-594.72,-61.486,-538.49,-64.303,-721.57
1951.000000000,8910.2,1297.5,1714.9,1643.0,1988.8,1068.5,2882.9,424.61,1601.2,288.75,648.35,740.12,0.0000,-3379.5,-6456.2,-274.13,-2530.5,-2351.1,-13462.,-1688.0,-1269.4,-5111.5,-2643.9,-5645.9,29870.,13351.,10227.,9598.8,18608.,6412.1,22984.,6641.8,10154.,3030.8,4355.7,5246.7,0.0000,-29.065,-30.327,-4.8357,-28.102,-16.736,-115.71,-93.559,-9.6714,-84.702,-10.114,-113.50
1952.000000000,8830.3,1290.8,1706.8,1638.8,1982.0,1055.3,2891.6,424.61,1587.9,289.49,645.81,744.78,0.0000,-3351.1,-6450.9,-272.45,-2530.2,-2330.8,-13461.,-1681.5,-1261.2,-5100.7,-2641.6,-5638.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1953.000000000,8815.9,1312.3,1709.4,1641.7,2001.9,1069.6,2908.0,429.59,1584.4,291.00,652.00,743.65,0.0000,-3344.3,-6442.2,-270.55,-2530.4,-2327.8,-13461.,-1676.5,-1256.7,-5096.3,-2641.1,-5635.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1954.000000000,8815.7,1299.6,1713.3,1640.6,1994.7,1057.6,2913.4,428.51,1580.5,290.54,656.38,744.64,0.0000,-3339.9,-6434.8,-269.06,-2530.3,-2325.5,-13462.,-1672.9,-1253.7,-5093.7,-2640.5,-5632.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1955.000000000,8809.4,1296.3,1722.0,1634.9,1985.2,1054.1,2911.6,427.24,1580.8,293.06,656.79,745.77,0.0000,-3335.9,-6427.5,-267.96,-2530.0,-2323.4,-13462.,-1670.3,-1251.4,-5092.2,-2640.1,-5630.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1956.000000000,8797.9,1280.5,1715.0,1644.5,1984.9,1050.3,2903.2,423.11,1578.8,292.11,653.60,746.64,0.0000,-3331.9,-6420.7,-267.15,-2529.5,-2321.2,-13461.,-1668.5,-1249.4,-5090.8,-2639.6,-5628.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1957.000000000,8801.1,1274.6,1702.0,1641.8,1949.1,1045.2,2884.6,419.61,1578.1,292.17,655.31,751.28,0.0000,-3328.0,-6414.3,-266.53,-2529.2,-2318.9,-13460.,-1667.2,-1247.6,-5089.6,-2639.4,-5626.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1958.000000000,8797.6,1273.9,1691.7,1624.9,1954.3,1050.3,2889.4,418.20,1576.8,292.25,654.44,749.95,0.0000,-3324.5,-6408.4,-266.03,-2529.0,-2316.7,-13459.,-1666.3,-1246.1,-5088.6,-2639.1,-5625.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1959.000000000,8784.7,1271.4,1695.9,1627.1,1943.2,1041.2,2885.5,415.61,1572.2,291.71,652.43,749.80,0.0000,-3321.1,-6403.2,-265.62,-2528.7,-2314.5,-13458.,-1665.7,-1244.8,-5087.6,-2638.6,-5624.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1960.000000000,8786.0,1262.5,1688.2,1623.6,1946.2,1039.0,2887.3,417.22,1575.0,292.55,652.18,749.24,0.0000,-3317.5,-6398.2,-265.27,-2528.2,-2312.3,-13456.,-1665.2,-1243.6,-5086.7,-2637.9,-5623.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1961.000000000,8777.1,1268.7,1676.3,1634.8,1945.4,1035.3,2894.4,419.55,1565.7,291.68,651.76,744.19,0.0000,-3314.2,-6393.9,-264.96,-2527.7,-2310.3,-13455.,-1664.8,-1242.5,-5085.9,-2637.6,-5622.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1962.000000000,8770.6,1262.1,1685.1,1638.7,1931.4,1035.2,2900.8,421.18,1548.8,288.76,651.95,746.11,0.0000,-3311.1,-6390.4,-264.69,-2527.2,-2308.4,-13454.,-1664.6,-1241.5,-5085.2,-2637.3,-5621.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1963.000000000,8771.9,1262.4,1688.6,1642.3,1936.3,1032.2,2885.9,422.08,1548.3,289.59,650.47,750.63,0.0000,-3308.1,-6387.5,-264.45,-2526.6,-2306.6,-13453.,-1664.3,-1240.7,-5084.7,-2637.0,-5621.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1964.000000000,8770.1,1258.9,1691.2,1651.8,1937.8,1038.7,2880.6,420.78,1549.1,291.79,650.94,749.05,0.0000,-3346.6,-6407.6,-268.15,-2526.1,-2332.0,-13452.,-1664.4,-1250.4,-5095.6,-2639.1,-5628.4,1410.8,630.58,483.05,453.35,878.85,302.85,1085.5,313.69,479.56,143.14,205.72,247.80,0.0000,-1.3683,-1.4294,-0.22839,-1.3257,-0.78808,-5.4644,-4.4208,-0.45678,-4.0009,-0.47765,-5.3646
1965.000000000,8774.9,1242.2,1658.7,1651.2,1938.0,1026.2,2879.8,417.53,1535.0,290.40,648.63,751.17,0.0000,-3322.8,-6406.7,-267.81,-2525.5,-2313.6,-13451.,-1664.3,-1246.7,-5087.3,-2637.5,-5622.7,77.618,34.694,26.576,24.943,48.352,16.662,59.724,17.259,26.385,7.8755,11.318,13.634,0.0000,-0.75270E-01,-0.78642E-01,-0.12566E-01,-0.72932E-01,-0.43287E-01,-0.30060,-0.24321,-0.25131E-01,-0.22012,-0.26278E-01,-0.29514
1966.000000000,8749.9,1255.5,1653.4,1656.3,1943.1,1035.3,2869.2,417.89,1562.4,290.17,645.69,749.01,0.0000,-3358.1,-6425.2,-270.83,-2525.1,-2336.8,-13450.,-1666.5,-1256.8,-5096.7,-2639.4,-5629.3,17524.,7832.8,6000.1,5631.3,10916.,3761.8,13484.,3896.5,5956.8,1778.0,2555.4,3078.1,0.0000,-17.017,-17.764,-2.8369,-16.477,-9.7889,-67.859,-54.907,-5.6739,-49.695,-5.9329,-66.631
1967.000000000,8656.3,1254.1,1688.4,1671.8,1863.2,1043.4,2864.2,420.75,1550.1,290.13,646.85,748.97,0.0000,-3374.7,-6445.6,-273.81,-2524.9,-2345.1,-13449.,-1690.0,-1265.5,-5104.4,-2640.2,-5638.0,0.18211E+06,81401.,62355.,58522.,0.11345E+06,39094.,0.14013E+06,40494.,61906.,18478.,26556.,31988.,0.0000,-177.15,-184.74,-29.482,-171.37,-101.85,-705.14,-570.71,-58.965,-516.45,-61.656,-692.46
1968.000000000,8657.9,1248.4,1687.4,1683.0,1810.9,1043.1,2859.5,422.51,1543.7,285.98,648.19,751.36,0.0000,-3388.6,-6463.9,-276.24,-2524.7,-2351.5,-13449.,-1683.9,-1273.3,-5107.5,-2640.7,-5642.1,4180.1,1868.4,1431.3,1343.3,2604.0,897.34,3216.5,929.48,1421.0,424.14,609.56,734.25,0.0000,-4.0743,-4.2443,-0.67672,-3.9369,-2.3399,-16.186,-13.101,-1.3534,-11.855,-1.4152,-15.895
1969.000000000,8638.5,1257.1,1695.1,1681.4,1933.9,1049.2,2890.8,428.48,1530.1,289.09,644.19,761.99,0.0000,-3359.8,-6457.3,-274.28,-2525.0,-2331.3,-13447.,-1678.3,-1264.1,-5096.3,-2638.7,-5634.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1970.000000000,8672.2,1290.6,1696.7,1676.7,1972.9,1055.1,2903.3,427.75,1516.9,288.91,644.03,761.92,0.0000,-3352.9,-6448.4,-272.17,-2525.2,-2327.6,-13448.,-1674.1,-1259.2,-5091.8,-2638.0,-5631.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1971.000000000,8693.0,1290.4,1705.5,1674.2,1970.5,1034.2,2903.2,421.96,1514.4,292.27,648.21,761.28,0.0000,-3348.2,-6439.8,-270.53,-2525.1,-2324.8,-13448.,-1671.0,-1255.8,-5089.7,-2637.4,-5628.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1972.000000000,8771.7,1278.8,1703.2,1674.1,1960.8,1021.4,2892.8,422.30,1516.3,294.58,640.07,760.42,0.0000,-3343.1,-6430.8,-269.31,-2524.8,-2321.9,-13447.,-1668.7,-1253.2,-5088.2,-2636.7,-5626.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1973.000000000,8795.7,1295.1,1571.7,1681.2,1959.9,1022.5,2906.1,425.51,1511.4,294.49,639.32,765.66,0.0000,-3339.2,-6422.9,-268.39,-2525.0,-2319.4,-13446.,-1667.2,-1251.1,-5086.7,-2636.7,-5624.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1974.000000000,8783.0,1304.2,1545.8,1681.8,1953.5,1029.2,2885.5,427.51,1514.9,292.83,642.68,770.50,0.0000,-3335.2,-6416.1,-267.70,-2524.7,-2317.2,-13446.,-1666.1,-1249.3,-5085.4,-2636.2,-5623.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1975.000000000,8787.5,1300.1,1555.2,1672.0,1951.0,1017.2,2852.9,428.25,1526.2,293.80,644.63,768.28,0.0000,-3331.4,-6411.3,-267.17,-2524.2,-2314.8,-13446.,-1665.4,-1247.7,-5084.6,-2636.1,-5622.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1976.000000000,8791.7,1298.0,1561.8,1669.1,1949.8,1009.0,2815.1,428.37,1528.5,295.29,645.73,766.14,0.0000,-3327.6,-6406.3,-266.74,-2523.6,-2312.4,-13445.,-1664.8,-1246.4,-5083.9,-2635.8,-5621.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1977.000000000,8790.8,1298.1,1565.1,1672.4,1951.1,1007.9,2801.8,425.26,1500.0,295.78,644.66,763.68,0.0000,-3323.8,-6401.6,-266.37,-2523.1,-2310.1,-13444.,-1664.4,-1245.1,-5083.1,-2635.9,-5620.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1978.000000000,8762.9,1298.9,1551.7,1672.4,1943.2,1008.4,2790.0,425.91,1497.8,292.87,640.63,763.03,0.0000,-3320.4,-6397.4,-266.04,-2522.6,-2308.0,-13443.,-1664.1,-1244.0,-5082.2,-2635.8,-5619.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1979.000000000,8757.7,1308.3,1538.2,1670.3,1949.5,1011.3,2801.9,423.26,1486.8,291.97,638.41,763.31,0.0000,-3317.5,-6393.5,-265.74,-2522.1,-2305.9,-13442.,-1663.9,-1243.0,-5081.4,-2635.6,-5619.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1980.000000000,8752.2,1306.8,1552.6,1670.6,1953.2,1007.1,2809.3,421.92,1484.7,292.62,636.49,760.78,0.0000,-3314.7,-6389.9,-265.47,-2521.6,-2304.0,-13441.,-1663.7,-1242.1,-5080.8,-2635.2,-5618.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1981.000000000,8735.2,1316.8,1583.1,1671.6,1992.1,1010.0,2824.7,423.69,1492.5,292.61,634.35,761.96,0.0000,-3353.3,-6409.6,-269.13,-2521.1,-2329.4,-13441.,-1664.9,-1252.1,-5091.8,-2637.2,-5626.3,9565.5,4275.6,3275.2,3073.9,5958.9,2053.4,7360.3,2126.9,3251.6,970.56,1394.9,1680.2,0.0000,-9.2842,-9.6913,-1.5486,-8.9947,-5.3246,-37.016,-29.984,-3.0971,-27.128,-3.2378,-36.389
1982.000000000,8742.9,1298.3,1627.1,1662.6,2074.8,997.55,2826.5,428.62,1487.5,291.45,629.99,761.17,0.0000,-3329.6,-6408.5,-268.74,-2520.6,-2311.0,-13441.,-1664.4,-1248.2,-5083.5,-2635.5,-5620.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1983.000000000,8743.2,1283.2,1630.0,1655.1,2074.2,995.12,2832.5,432.33,1481.0,291.22,625.29,760.26,0.0000,-3323.3,-6403.9,-267.81,-2520.1,-2307.0,-13440.,-1664.0,-1246.0,-5081.1,-2634.7,-5619.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1984.000000000,8712.1,1282.6,1631.0,1661.4,2078.8,1004.4,2844.7,434.21,1473.7,292.90,624.00,760.67,0.0000,-3319.3,-6399.0,-266.99,-2519.7,-2304.4,-13439.,-1663.7,-1244.4,-5079.9,-2633.9,-5618.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1985.000000000,8717.7,1291.2,1633.8,1646.6,2064.1,1006.3,2839.1,433.95,1470.5,293.73,621.20,759.73,0.0000,-3315.9,-6394.1,-266.32,-2519.3,-2302.2,-13439.,-1663.5,-1243.1,-5079.1,-2633.1,-5617.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1986.000000000,8721.1,1287.8,1629.9,1631.3,2041.3,1005.6,2838.1,434.65,1470.5,292.60,620.56,753.49,0.0000,-3312.8,-6389.7,-265.78,-2518.9,-2300.2,-13438.,-1663.3,-1242.0,-5078.4,-2632.3,-5617.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1987.000000000,8704.2,1282.5,1628.6,1635.3,2054.4,1006.5,2836.6,430.65,1474.1,291.77,620.54,752.89,0.0000,-3309.8,-6385.9,-265.33,-2518.6,-2298.3,-13438.,-1663.1,-1241.0,-5077.9,-2631.6,-5616.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1988.000000000,8628.7,1263.6,1617.7,1645.8,2086.9,1006.0,2827.4,428.65,1476.4,291.32,616.62,754.69,0.0000,-3306.8,-6382.0,-264.94,-2518.3,-2296.3,-13438.,-1663.1,-1240.2,-5077.4,-2630.6,-5616.6,400.01,178.80,136.96,128.54,249.19,85.868,307.79,88.944,135.97,40.587,58.330,70.262,0.0000,-0.38695,-0.40467,-0.64758E-01,-0.37555,-0.22142,-1.5468,-1.2532,-0.12952,-1.1343,-0.13533,-1.5212
1989.000000000,8630.5,1267.0,1597.2,1642.0,2104.8,1003.3,2831.2,427.34,1468.6,291.62,616.53,760.29,0.0000,-3304.0,-6378.5,-264.60,-2518.0,-2294.4,-13437.,-1662.9,-1239.4,-5076.9,-2630.0,-5616.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1990.000000000,8519.6,1264.6,1613.2,1645.0,2085.3,1003.7,2831.8,428.52,1470.0,293.10,615.39,761.64,0.0000,-3301.0,-6375.7,-264.31,-2517.8,-2292.7,-13436.,-1662.8,-1238.6,-5076.6,-2629.6,-5616.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1991.000000000,8558.7,1268.8,1628.5,1645.9,2067.1,1000.4,2822.0,427.25,1475.4,295.81,614.15,765.81,0.0000,-3298.1,-6373.4,-264.04,-2517.6,-2291.0,-13435.,-1662.7,-1238.0,-5076.5,-2629.2,-5615.9,49.153,21.971,16.830,15.796,30.620,10.552,37.822,10.930,16.709,4.9874,7.1677,8.6339,0.0000,-0.47469E-01,-0.49686E-01,-0.79575E-02,-0.46115E-01,-0.27173E-01,-0.19001,-0.15396,-0.15915E-01,-0.13937,-0.16627E-01,-0.18691
1992.000000000,8589.5,1283.2,1638.1,1643.8,2048.7,1005.3,2797.9,425.35,1470.6,293.72,614.39,767.68,0.0000,-3295.2,-6371.5,-263.78,-2517.4,-2289.4,-13435.,-1662.6,-1237.4,-5076.3,-2628.9,-5615.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1993.000000000,8702.3,1286.6,1636.6,1653.0,2048.0,1011.4,2779.1,426.64,1472.8,293.59,612.59,769.45,0.0000,-3292.4,-6369.6,-263.52,-2517.1,-2287.8,-13434.,-1662.6,-1237.1,-5076.0,-2628.5,-5615.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1994.000000000,8708.1,1288.2,1643.0,1652.1,2039.7,1011.5,2807.9,427.32,1462.6,294.52,612.51,769.20,0.0000,-3289.9,-6367.7,-263.27,-2516.9,-2286.2,-13433.,-1662.5,-1236.8,-5075.7,-2628.1,-5615.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1995.000000000,8679.3,1286.1,1645.1,1658.0,2027.4,1006.4,2820.4,421.04,1458.5,292.69,614.74,768.84,0.0000,-3287.6,-6365.8,-263.02,-2516.7,-2284.7,-13432.,-1662.5,-1236.5,-5075.2,-2627.7,-5615.0,730.43,326.49,250.10,234.73,455.03,156.80,562.04,162.42,248.30,74.113,106.51,128.30,0.0000,-0.70386,-0.73759,-0.11825,-0.68471,-0.40323,-2.8229,-2.2872,-0.23650,-2.0710,-0.24704,-2.7770
1996.000000000,8773.8,1279.5,1652.8,1665.1,2017.3,1012.1,2843.2,421.53,1458.7,291.06,615.61,769.58,0.0000,-3326.8,-6386.9,-266.67,-2516.6,-2310.3,-13432.,-1664.2,-1244.5,-5086.6,-2629.8,-5623.1,12555.,5611.7,4298.7,4034.5,7821.0,2695.1,9660.4,2791.6,4267.7,1273.9,1830.8,2205.2,0.0000,-12.116,-12.683,-2.0325,-11.777,-6.9483,-48.517,-39.311,-4.0650,-35.595,-4.2462,-47.729
1997.000000000,8741.1,1254.1,1645.7,1654.4,2029.0,1004.8,2852.7,418.53,1449.2,290.13,618.11,767.72,0.0000,-3303.5,-6386.9,-266.28,-2516.6,-2292.3,-13431.,-1663.7,-1241.8,-5079.0,-2628.1,-5617.8,9.7928,4.3772,3.3530,3.1469,6.1005,2.1022,7.5352,2.1775,3.3289,0.99363,1.4280,1.7201,0.0000,-0.94508E-02,-0.98934E-02,-0.15854E-02,-0.91857E-02,-0.54135E-02,-0.37842E-01,-0.30661E-01,-0.31707E-02,-0.27764E-01,-0.33119E-02,-0.37227E-01
1998.000000000,8670.1,1244.5,1636.7,1645.5,2035.2,1003.2,2840.0,420.95,1457.8,288.92,617.84,765.54,0.0000,-3297.4,-6383.2,-265.35,-2516.4,-2288.7,-13431.,-1663.2,-1240.3,-5076.9,-2627.4,-5615.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
1999.000000000,8662.3,1252.9,1639.1,1647.2,2049.8,1013.3,2840.5,421.40,1468.0,288.85,618.62,764.82,0.0000,-3335.1,-6402.0,-268.42,-2516.7,-2313.8,-13431.,-1663.3,-1249.1,-5087.5,-2629.3,-5622.9,2511.8,1122.7,860.04,807.18,1564.8,539.21,1932.8,558.52,853.84,254.86,366.28,441.20,0.0000,-2.4267,-2.5386,-0.40664,-2.3575,-1.3905,-9.7050,-7.8632,-0.81328,-7.1212,-0.84947,-9.5480
2000.000000000,8659.1,1258.2,1624.0,1642.4,1962.5,999.58,2831.3,422.98,1457.3,288.86,614.49,763.14,0.0000,-3311.0,-6400.1,-267.60,-2517.0,-2295.6,-13430.,-1662.9,-1245.3,-5079.0,-2627.5,-5617.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
2001.000000000,8641.1,1261.6,1625.2,1640.1,1971.9,1001.7,2836.7,426.63,1453.2,288.88,610.53,767.22,0.0000,-3304.8,-6394.9,-266.37,-2517.1,-2291.7,-13429.,-1662.6,-1243.1,-5076.3,-2626.7,-5615.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
2002.000000000,8636.2,1252.5,1620.1,1634.7,1961.3,1007.4,2830.5,427.08,1467.9,287.80,606.35,766.70,0.0000,-3300.9,-6390.3,-265.34,-2517.1,-2289.5,-13428.,-1662.4,-1241.5,-5075.1,-2625.8,-5614.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
2003.000000000,8635.9,1252.0,1621.9,1627.7,1957.8,1006.0,2842.4,429.83,1478.1,288.81,606.81,762.65,0.0000,-3297.8,-6386.1,-264.54,-2516.9,-2287.7,-13427.,-1662.2,-1240.2,-5074.4,-2624.9,-5613.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
2004.000000000,8759.1,1262.8,1624.0,1632.8,1956.8,995.10,2839.8,432.78,1479.5,287.97,607.70,757.48,0.0000,-3294.9,-6381.7,-263.90,-2516.7,-2285.9,-13426.,-1662.1,-1239.2,-5073.5,-2624.1,-5612.5,191.15,85.442,65.451,61.428,119.08,41.034,147.09,42.504,64.979,19.395,27.875,33.576,0.0000,-0.18440,-0.19306,-0.30946E-01,-0.17925,-0.10537,-0.73832,-0.59818,-0.61892E-01,-0.54186,-0.64632E-01,-0.72645
2005.000000000,8716.7,1270.1,1626.2,1635.2,1960.4,986.50,2820.2,427.63,1476.2,286.51,608.34,755.36,0.0000,-3292.3,-6377.6,-263.40,-2516.7,-2284.2,-13425.,-1662.0,-1238.2,-5072.8,-2623.3,-5611.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
2006.000000000,8544.3,1265.9,1626.0,1637.3,1964.7,993.49,2809.6,422.95,1481.4,284.31,609.72,758.61,0.0000,-3289.7,-6374.1,-262.98,-2516.7,-2282.7,-13425.,-1661.9,-1237.2,-5072.2,-2622.7,-5611.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
2007.000000000,8461.6,1263.9,1617.4,1636.7,1974.4,1020.9,2810.8,424.82,1480.3,285.58,612.49,758.33,0.0000,-3328.5,-6393.7,-266.52,-2516.9,-2308.6,-13425.,-1663.2,-1245.4,-5083.4,-2624.7,-5619.0,10567.,4723.3,3618.2,3395.8,6582.9,2268.4,8131.1,2349.7,3592.1,1072.2,1540.9,1856.1,0.0000,-10.198,-10.670,-1.7107,-9.9113,-5.8330,-40.804,-33.061,-3.4214,-29.953,-3.5727,-40.154
2008.000000000,8471.6,1256.2,1597.3,1648.0,1969.7,1019.3,2798.4,425.88,1478.6,284.76,613.98,760.95,0.0000,-3304.9,-6392.6,-266.06,-2516.9,-2290.7,-13424.,-1662.8,-1242.0,-5075.2,-2623.0,-5613.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
2009.000000000,8466.0,1250.9,1590.3,1652.7,1938.0,1021.8,2794.7,430.09,1494.7,282.01,610.63,761.23,0.0000,-3298.7,-6387.9,-265.08,-2516.9,-2287.1,-13423.,-1662.4,-1240.1,-5072.5,-2622.3,-5611.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
2010.000000000,8465.3,1255.5,1589.0,1648.5,1875.5,1016.7,2804.7,433.93,1504.2,278.82,605.40,761.59,0.0000,-3294.9,-6382.8,-264.22,-2516.7,-2284.9,-13422.,-1662.1,-1238.7,-5071.1,-2621.7,-5610.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
2011.000000000,8463.5,1259.6,1596.3,1652.0,1855.5,1021.3,2820.9,433.62,1503.0,278.34,601.66,760.88,0.0000,-3291.5,-6378.1,-263.54,-2516.2,-2283.0,-13421.,-1661.9,-1237.6,-5070.2,-2621.2,-5610.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
2012.000000000,8470.8,1260.4,1607.3,1653.5,1858.1,1038.5,2816.0,433.46,1504.5,276.35,604.51,760.92,0.0000,-3329.9,-6396.7,-266.90,-2515.8,-2308.5,-13421.,-1664.3,-1246.1,-5081.5,-2623.1,-5618.1,19148.,8558.9,6556.3,6153.3,11928.,4110.5,14734.,4257.7,6509.1,1942.9,2792.3,3363.4,0.0000,-18.482,-19.330,-3.0999,-17.962,-10.562,-73.904,-59.888,-6.1998,-54.271,-6.4731,-72.747
2013.000000000,8437.4,1255.2,1604.1,1651.8,1836.4,1039.7,2801.3,433.46,1502.1,273.88,603.39,758.25,0.0000,-3347.4,-6417.3,-270.23,-2515.6,-2317.6,-13421.,-1668.0,-1254.4,-5085.6,-2623.8,-5621.9,33279.,14875.,11395.,10694.,20731.,7143.8,25607.,7399.7,11312.,3376.6,4852.8,5845.4,0.0000,-32.178,-33.618,-5.3875,-31.242,-18.387,-128.43,-104.08,-10.775,-94.319,-11.250,-126.43
2014.000000000,8406.3,1257.2,1603.2,1651.3,1820.0,1044.0,2810.1,436.10,1514.6,274.49,598.95,753.66,0.0000,-3361.5,-6436.2,-272.93,-2515.5,-2324.5,-13421.,-1676.6,-1262.0,-5089.3,-2624.1,-5626.2,77706.,34733.,26607.,24971.,48408.,16681.,59792.,17279.,26415.,7884.5,11331.,13649.,0.0000,-75.282,-78.566,-12.580,-73.013,-42.992,-299.86,-243.04,-25.160,-220.24,-26.269,-295.21
2015.000000000,8388.2,1263.0,1603.2,1659.2,1813.2,1045.5,2810.6,438.01,1513.4,274.22,600.17,754.77,0.0000,-3374.5,-6453.2,-275.07,-2515.5,-2330.7,-13420.,-1683.6,-1269.1,-5092.8,-2624.3,-5630.7,82060.,36679.,28097.,26370.,51120.,17616.,63143.,18247.,27895.,8326.3,11966.,14414.,0.0000,-79.660,-83.044,-13.285,-77.171,-45.453,-316.64,-256.69,-26.570,-232.58,-27.741,-311.76
2016.000000000,8380.6,1265.7,1602.5,1665.4,1810.9,1058.0,2818.3,440.28,1511.5,274.69,600.97,760.32,0.0000,-3386.8,-6468.5,-276.81,-2515.4,-2336.6,-13420.,-1682.3,-1275.7,-5094.6,-2624.3,-5633.3,34806.,15557.,11917.,11185.,21682.,7471.6,26782.,7739.3,11831.,3531.5,5075.5,6113.7,0.0000,-33.857,-35.259,-5.6347,-32.760,-19.299,-134.31,-108.89,-11.269,-98.649,-11.766,-132.24
2017.000000000,8367.2,1273.9,1601.1,1659.0,1818.3,1077.0,2854.9,442.69,1515.8,275.72,604.29,767.61,0.0000,-3399.0,-6482.1,-278.29,-2515.7,-2343.3,-13421.,-1684.2,-1281.9,-5096.1,-2624.5,-5635.3,57614.,25752.,19727.,18514.,35891.,12368.,44332.,12811.,19585.,5845.8,8401.4,10120.,0.0000,-56.185,-58.439,-9.3272,-54.305,-32.040,-222.42,-180.29,-18.654,-163.31,-19.478,-218.97
2018.000000000,8323.0,1289.4,1601.7,1632.0,1821.9,1054.8,2863.8,444.45,1505.7,273.48,610.44,759.41,0.0000,-3370.1,-6472.5,-275.66,-2516.1,-2322.8,-13421.,-1677.9,-1270.2,-5084.3,-2622.4,-5627.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
2019.000000000,8312.0,1268.8,1609.6,1621.2,1800.4,1045.1,2857.7,444.89,1496.2,276.45,622.62,763.86,0.0000,-3361.3,-6460.9,-273.08,-2516.4,-2318.4,-13422.,-1673.1,-1263.9,-5080.1,-2621.6,-5622.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
2020.000000000,8313.6,1268.8,1624.5,1618.6,1800.7,1041.9,2849.9,443.46,1499.3,278.92,627.95,760.56,0.0000,-3355.6,-6450.4,-271.10,-2516.4,-2315.8,-13423.,-1669.7,-1259.5,-5078.1,-2621.2,-5619.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
2021.000000000,8249.7,1250.0,1622.0,1611.1,1793.7,1026.9,2820.0,442.58,1509.7,278.62,625.07,756.23,0.0000,-3350.3,-6439.7,-269.64,-2516.6,-2312.7,-13423.,-1667.2,-1256.1,-5076.7,-2621.3,-5616.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
2022.000000000,8203.7,1253.4,1616.7,1612.3,1779.1,1009.7,2795.7,440.16,1508.7,275.08,624.07,759.41,0.0000,-3345.6,-6430.0,-268.54,-2516.9,-2309.7,-13422.,-1665.5,-1253.3,-5075.2,-2621.2,-5614.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
2023.000000000,8280.2,1243.5,1712.4,1612.7,1763.3,999.92,2781.2,439.82,1511.8,274.13,628.39,762.23,0.0000,-3340.4,-6421.0,-267.70,-2516.6,-2306.8,-13420.,-1664.3,-1250.9,-5074.0,-2620.7,-5613.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
2024.000000000,8281.6,1234.0,1703.3,1631.7,1753.8,1004.5,2789.9,440.76,1514.7,270.72,629.52,758.24,0.0000,-3335.8,-6413.9,-267.05,-2516.3,-2304.2,-13420.,-1663.4,-1248.9,-5072.9,-2620.9,-5612.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
2025.000000000,8222.3,1226.7,1694.8,1637.1,1766.5,1006.7,2799.2,441.43,1512.5,268.91,631.35,759.48,0.0000,-3331.4,-6408.0,-266.54,-2515.8,-2301.8,-13419.,-1662.8,-1247.1,-5072.2,-2620.9,-5610.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
2026.000000000,8228.6,1227.7,1693.8,1647.9,1764.4,1004.9,2814.3,439.47,1503.0,268.25,632.08,757.12,0.0000,-3327.1,-6402.5,-266.13,-2515.0,-2299.3,-13418.,-1662.4,-1245.5,-5071.6,-2621.0,-5609.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
2027.000000000,8200.6,1229.5,1699.3,1640.8,1763.8,1007.6,2815.1,442.61,1498.9,270.93,634.39,760.92,0.0000,-3322.9,-6397.9,-265.77,-2514.2,-2296.9,-13417.,-1662.0,-1244.1,-5071.0,-2621.5,-5609.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
2028.000000000,8056.6,1226.2,1694.9,1631.8,1756.3,997.31,2821.6,445.47,1494.1,272.28,636.98,760.79,0.0000,-3318.8,-6392.9,-265.44,-2513.5,-2294.6,-13416.,-1661.8,-1242.8,-5070.3,-2621.9,-5608.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
2029.000000000,8039.2,1220.2,1699.9,1630.9,1761.7,989.52,2825.1,446.35,1487.4,271.55,624.45,759.78,0.0000,-3315.6,-6387.7,-265.13,-2512.9,-2292.3,-13415.,-1661.6,-1241.5,-5069.4,-2621.6,-5608.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
2030.000000000,8056.8,1209.9,1700.0,1635.2,1790.6,983.13,2811.9,444.65,1486.0,269.68,618.23,749.71,0.0000,-3312.4,-6382.4,-264.84,-2512.3,-2290.0,-13414.,-1661.4,-1240.4,-5068.7,-2620.9,-5607.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
2031.000000000,8028.2,1199.9,1694.0,1634.9,1789.9,984.61,2809.9,445.70,1496.5,269.07,616.33,750.55,0.0000,-3309.2,-6377.9,-264.55,-2511.7,-2287.8,-13414.,-1661.3,-1239.4,-5068.1,-2620.3,-5607.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
2032.000000000,8129.5,1187.4,1689.9,1653.8,1794.5,982.02,2790.2,447.82,1502.1,268.30,617.14,750.09,0.0000,-3305.9,-6374.0,-264.28,-2511.0,-2285.8,-13413.,-1661.2,-1238.5,-5067.4,-2619.7,-5606.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
2033.000000000,8165.3,1187.1,1672.8,1662.2,1788.4,985.19,2794.4,448.71,1507.4,268.68,610.17,750.28,0.0000,-3302.7,-6370.6,-264.03,-2510.3,-2283.8,-13413.,-1661.1,-1237.7,-5066.9,-2619.2,-5606.4,0.46730,0.20888,0.16000,0.15017,0.29111,0.10031,0.35957,0.10391,0.15885,0.47415E-01,0.68144E-01,0.82082E-01,0.0000,-0.45188E-03,-0.47209E-03,-0.75652E-04,-0.43881E-03,-0.25733E-03,-0.18026E-02,-0.14629E-02,-0.15130E-03,-0.13246E-02,-0.15796E-03,-0.17770E-02
2034.000000000,8171.6,1199.6,1660.0,1665.6,1808.6,986.15,2802.3,448.46,1506.3,268.21,602.95,748.99,0.0000,-3299.8,-6367.4,-263.78,-2509.6,-2281.8,-13413.,-1661.0,-1236.9,-5066.4,-2618.8,-5606.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
2035.000000000,8187.2,1192.2,1658.5,1657.0,1779.9,984.78,2800.1,451.62,1499.6,269.96,600.81,746.64,0.0000,-3296.9,-6364.7,-263.53,-2508.9,-2279.9,-13412.,-1660.9,-1236.2,-5065.8,-2618.3,-5605.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
2036.000000000,8170.4,1198.7,1668.6,1650.1,1762.6,984.23,2809.7,455.46,1497.5,269.38,602.70,746.17,0.0000,-3294.2,-6362.2,-263.28,-2508.3,-2278.0,-13413.,-1660.8,-1235.5,-5065.3,-2617.8,-5605.7,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
2037.000000000,8163.3,1191.6,1671.4,1660.2,1759.2,982.44,2812.3,451.51,1480.3,269.87,601.51,746.87,0.0000,-3291.7,-6359.7,-263.02,-2507.7,-2276.1,-13413.,-1660.8,-1234.9,-5064.8,-2617.1,-5605.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
2038.000000000,8019.6,1197.6,1680.3,1659.8,1759.9,996.13,2805.4,450.36,1474.8,270.32,600.73,746.55,0.0000,-3330.6,-6380.3,-266.65,-2507.3,-2301.5,-13414.,-1685.6,-1243.1,-5080.9,-2619.0,-5619.7,0.18709E+06,83627.,64061.,60123.,0.11655E+06,40163.,0.14396E+06,41602.,63599.,18983.,27283.,32863.,0.0000,-180.75,-188.83,-30.289,-175.61,-103.01,-721.41,-585.64,-60.577,-530.27,-63.227,-711.35
2039.000000000,7983.5,1199.5,1682.7,1661.9,1759.2,1002.6,2781.9,453.06,1473.0,271.02,596.71,748.08,0.0000,-3348.8,-6403.0,-270.15,-2507.0,-2310.4,-13415.,-1680.1,-1251.2,-5086.7,-2619.5,-5625.7,5325.5,2380.4,1823.4,1711.4,3317.5,1143.2,4097.8,1184.2,1810.3,540.35,776.58,935.43,0.0000,-5.1543,-5.3785,-0.86215,-5.0026,-2.9369,-20.534,-16.671,-1.7243,-15.094,-1.7997,-20.249
2040.000000000,7994.3,1197.2,1661.8,1667.5,1752.4,997.49,2783.4,450.14,1473.6,269.58,591.11,746.18,0.0000,-3321.9,-6400.7,-269.04,-2506.8,-2289.9,-13415.,-1674.7,-1246.2,-5076.3,-2617.0,-5619.0,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
2041.000000000,7940.7,1209.1,1651.4,1675.1,1764.1,1016.1,2805.3,449.58,1464.8,268.55,589.70,748.54,0.0000,-3315.0,-6394.3,-267.49,-2506.9,-2286.5,-13415.,-1670.6,-1243.5,-5072.3,-2616.2,-5615.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
2042.000000000,7848.3,1223.6,1643.7,1671.4,1778.4,1011.8,2814.0,450.13,1465.4,268.92,593.89,742.99,0.0000,-3311.3,-6389.1,-266.22,-2506.9,-2284.3,-13416.,-1667.6,-1241.7,-5070.0,-2615.9,-5613.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
2043.000000000,7968.9,1207.1,1641.2,1663.1,1894.0,1008.0,2810.3,448.24,1456.3,273.23,592.30,745.81,0.0000,-3307.5,-6383.6,-265.25,-2506.7,-2282.2,-13416.,-1665.5,-1240.2,-5068.9,-2615.7,-5611.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
2044.000000000,7989.5,1204.0,1636.5,1660.2,1905.0,1007.5,2809.3,448.41,1454.6,273.49,592.39,745.26,0.0000,-3303.9,-6379.0,-264.50,-2506.4,-2280.3,-13415.,-1664.1,-1239.0,-5067.9,-2615.5,-5609.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
2045.000000000,7969.6,1192.2,1643.4,1660.1,1904.8,1003.6,2769.7,448.55,1451.9,273.27,592.43,744.58,0.0000,-3300.8,-6374.9,-263.90,-2506.3,-2278.3,-13414.,-1663.0,-1238.0,-5067.2,-2615.6,-5608.3,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
2046.000000000,7959.0,1198.1,1640.3,1665.3,1909.9,1003.7,2762.5,449.80,1446.9,273.64,597.05,751.47,0.0000,-3297.4,-6371.2,-263.40,-2506.1,-2276.0,-13413.,-1662.3,-1237.2,-5066.5,-2615.2,-5607.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
2047.000000000,7932.9,1199.2,1652.9,1655.6,1905.4,1008.4,2750.5,451.14,1442.1,273.67,598.86,750.81,0.0000,-3294.1,-6367.0,-262.97,-2505.8,-2274.0,-13411.,-1661.8,-1236.5,-5065.8,-2614.9,-5606.6,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
2048.000000000,7916.1,1193.9,1648.0,1644.4,1897.2,1007.5,2757.5,447.56,1435.4,270.82,597.72,747.55,0.0000,-3291.1,-6363.5,-262.59,-2505.5,-2272.2,-13410.,-1661.5,-1235.8,-5065.0,-2614.8,-5606.0,839.33,375.16,287.39,269.72,522.87,180.18,645.84,186.63,285.31,85.163,122.39,147.43,0.0000,-0.80969,-0.84634,-0.13588,-0.78716,-0.46110,-3.2362,-2.6279,-0.27176,-2.3789,-0.28358,-3.1924
2049.000000000,7906.7,1190.6,1639.8,1649.5,1894.5,1014.5,2750.9,447.48,1438.3,270.33,602.93,746.17,0.0000,-3329.9,-6383.8,-266.17,-2505.3,-2297.7,-13410.,-1670.7,-1244.1,-5077.9,-2617.3,-5615.8,71030.,31749.,24320.,22826.,44248.,15248.,54655.,15794.,24145.,7207.0,10358.,12476.,0.0000,-68.612,-71.648,-11.499,-66.657,-39.108,-273.85,-222.40,-22.998,-201.31,-24.000,-270.16
2050.000000000,7903.6,1193.6,1649.2,1647.4,1892.6,1021.6,2726.1,450.55,1438.4,270.54,605.17,745.98,0.0000,-3347.6,-6405.8,-269.65,-2505.1,-2306.7,-13410.,-1674.8,-1252.1,-5083.5,-2618.2,-5621.0,49419.,22089.,16921.,15881.,30786.,10609.,38027.,10989.,16799.,5014.3,7206.5,8680.6,0.0000,-47.822,-49.884,-8.0005,-46.414,-27.251,-190.52,-154.74,-16.001,-140.07,-16.699,-187.96
2051.000000000,7914.2,1201.1,1651.6,1669.5,1895.5,1024.4,2719.1,450.39,1444.8,269.95,610.26,746.40,0.0000,-3361.9,-6426.3,-272.47,-2505.0,-2313.8,-13410.,-1679.7,-1259.8,-5087.1,-2619.1,-5625.0,65417.,29240.,22399.,21022.,40752.,14043.,50336.,14546.,22237.,6637.5,9539.3,11491.,0.0000,-63.424,-66.087,-10.590,-61.492,-36.116,-252.18,-204.85,-21.181,-185.41,-22.105,-248.81
2052.000000000,7900.6,1187.6,1654.6,1673.2,1909.3,1031.9,2721.5,453.53,1447.2,270.46,613.02,748.16,0.0000,-3375.2,-6445.1,-274.70,-2505.5,-2320.1,-13409.,-1676.7,-1266.9,-5088.5,-2620.1,-5626.7,15773.,7050.3,5400.7,5068.8,9826.0,3386.0,12137.,3507.3,5361.8,1600.4,2300.1,2770.6,0.0000,-15.323,-15.950,-2.5535,-14.839,-8.7167,-60.807,-49.396,-5.1071,-44.705,-5.3300,-59.996
2053.000000000,7836.4,1183.8,1644.0,1665.9,1915.1,1030.6,2764.6,457.94,1432.8,273.40,611.77,758.25,0.0000,-3346.4,-6438.5,-272.58,-2506.3,-2299.7,-13409.,-1672.2,-1258.1,-5076.7,-2618.3,-5618.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
2054.000000000,7891.4,1217.2,1648.2,1660.5,1922.0,1050.0,2780.8,459.34,1425.8,272.02,615.54,756.44,0.0000,-3339.7,-6429.6,-270.34,-2507.1,-2296.2,-13410.,-1668.8,-1253.3,-5072.3,-2618.0,-5614.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
2055.000000000,7894.4,1194.3,1649.0,1656.1,1919.6,1045.4,2764.4,453.32,1421.0,273.03,615.51,755.45,0.0000,-3335.0,-6420.7,-268.59,-2507.4,-2293.4,-13411.,-1666.4,-1250.0,-5070.4,-2617.3,-5611.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
2056.000000000,7893.1,1208.7,1629.5,1656.9,1941.4,1032.5,2755.2,451.55,1408.1,273.35,611.86,752.67,0.0000,-3330.8,-6411.9,-267.27,-2507.7,-2290.6,-13411.,-1664.6,-1247.4,-5068.7,-2616.6,-5609.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
2057.000000000,8001.4,1210.6,1631.1,1660.9,1950.4,1019.2,2733.3,447.79,1409.8,271.63,609.49,750.22,0.0000,-3326.9,-6403.2,-266.28,-2508.2,-2287.9,-13411.,-1663.4,-1245.3,-5067.2,-2615.7,-5608.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
2058.000000000,8012.5,1227.2,1626.5,1653.3,1954.4,1037.2,2725.1,449.49,1418.2,273.96,607.77,750.34,0.0000,-3364.8,-6418.5,-269.43,-2508.6,-2312.8,-13412.,-1664.7,-1255.8,-5077.9,-2617.3,-5615.2,15532.,6942.4,5318.0,4991.2,9675.6,3334.1,11951.,3453.6,5279.7,1575.9,2264.9,2728.2,0.0000,-15.095,-15.712,-2.5144,-14.616,-8.5892,-59.912,-48.663,-5.0289,-44.024,-5.2485,-59.110
2059.000000000,8017.3,1238.8,1624.5,1664.2,1953.6,1042.4,2738.7,447.80,1420.8,272.70,611.98,746.53,0.0000,-3381.9,-6437.5,-272.61,-2509.0,-2321.4,-13413.,-1667.6,-1264.3,-5081.9,-2618.3,-5618.2,29840.,13338.,10217.,9589.1,18589.,6405.6,22961.,6635.1,10143.,3027.7,4351.3,5241.4,0.0000,-29.049,-30.204,-4.8308,-28.101,-16.524,-115.09,-93.494,-9.6615,-84.579,-10.084,-113.56
2060.000000000,8082.3,1230.4,1623.9,1660.4,1955.6,1027.5,2730.7,446.33,1408.5,269.97,618.48,743.83,0.0000,-3353.8,-6432.7,-271.29,-2509.1,-2300.4,-13413.,-1665.7,-1256.5,-5071.8,-2616.5,-5611.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
2061.000000000,8226.3,1225.2,1628.4,1663.8,1944.4,1025.5,2698.1,448.09,1401.1,272.42,621.30,742.48,0.0000,-3345.1,-6424.2,-269.60,-2508.9,-2295.4,-13412.,-1664.2,-1252.1,-5068.6,-2616.1,-5608.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
2062.000000000,8278.5,1224.7,1646.5,1668.8,1947.2,1027.5,2672.7,452.16,1398.5,271.99,623.95,744.37,0.0000,-3339.2,-6415.9,-268.23,-2508.5,-2292.2,-13412.,-1663.1,-1249.1,-5067.0,-2616.1,-5607.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
2063.000000000,8254.4,1234.0,1647.4,1669.1,1944.4,1028.8,2671.2,446.91,1393.3,268.17,611.60,746.06,0.0000,-3334.4,-6408.7,-267.18,-2508.2,-2289.6,-13411.,-1662.3,-1246.7,-5065.3,-2615.8,-5606.1,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
2064.000000000,8250.3,1233.9,1651.1,1685.5,1944.2,1033.9,2674.7,445.54,1390.3,266.26,611.75,740.17,0.0000,-3330.0,-6401.9,-266.36,-2507.8,-2287.0,-13410.,-1661.7,-1244.6,-5064.1,-2615.3,-5605.2,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
2065.000000000,8229.6,1221.5,1646.4,1685.2,1939.7,1048.3,2683.9,446.93,1388.5,266.01,612.86,738.38,0.0000,-3325.5,-6395.4,-265.72,-2507.3,-2284.6,-13410.,-1661.3,-1242.9,-5063.1,-2615.1,-5604.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
2066.000000000,8183.8,1202.1,1654.2,1680.9,1948.2,1054.9,2712.0,449.42,1399.9,266.50,610.68,740.75,0.0000,-3321.2,-6389.8,-265.18,-2506.9,-2282.5,-13410.,-1661.0,-1241.4,-5062.5,-2614.9,-5603.8,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
2067.000000000,8170.2,1203.9,1651.3,1673.2,1942.3,1049.0,2716.3,450.86,1408.3,267.38,609.14,741.89,0.0000,-3317.2,-6384.9,-264.73,-2506.5,-2280.6,-13409.,-1660.7,-1240.1,-5062.1,-2614.8,-5603.4,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
2068.000000000,8154.7,1203.5,1639.3,1670.5,1933.7,1052.4,2725.2,452.89,1407.8,266.60,603.96,745.05,0.0000,-3313.6,-6380.5,-264.33,-2506.1,-2278.7,-13409.,-1660.6,-1239.3,-5061.6,-2614.4,-5602.9,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
2069.000000000,8155.5,1184.9,1646.8,1663.7,1930.9,1049.1,2734.3,448.86,1410.9,264.90,597.91,742.96,0.0000,-3310.6,-6376.7,-263.97,-2505.8,-2276.8,-13409.,-1660.4,-1238.5,-5060.9,-2613.7,-5602.5,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000,0.0000
