time,RECHARGE
1.000000000000,0.0000
2.000000000000,0.0000
3.000000000000,0.0000
4.000000000000,759.37
5.000000000000,400.14
6.000000000000,0.0000
7.000000000000,0.0000
8.000000000000,10.434
9.000000000000,4519.5
10.00000000000,5266.5
11.00000000000,0.0000
12.00000000000,0.0000
13.00000000000,0.0000
14.00000000000,0.0000
15.00000000000,0.0000
16.00000000000,0.0000
17.00000000000,0.0000
18.00000000000,0.0000
19.00000000000,0.0000
20.00000000000,0.0000
21.00000000000,0.0000
22.00000000000,0.0000
23.00000000000,0.0000
24.00000000000,0.0000
25.00000000000,0.0000
26.00000000000,0.0000
27.00000000000,0.0000
28.00000000000,0.0000
29.00000000000,0.0000
30.00000000000,0.0000
31.00000000000,0.0000
32.00000000000,0.0000
33.00000000000,0.0000
34.00000000000,0.0000
35.00000000000,0.0000
36.00000000000,0.0000
37.00000000000,0.0000
38.00000000000,0.0000
39.00000000000,0.0000
40.00000000000,0.0000
41.00000000000,29.940
42.00000000000,0.0000
43.00000000000,0.0000
44.00000000000,0.0000
45.00000000000,0.0000
46.00000000000,0.0000
47.00000000000,0.0000
48.00000000000,0.0000
49.00000000000,0.0000
50.00000000000,0.0000
51.00000000000,0.0000
52.00000000000,257.46
53.00000000000,0.0000
54.00000000000,0.0000
55.00000000000,0.0000
56.00000000000,248.88
57.00000000000,0.0000
58.00000000000,0.0000
59.00000000000,0.0000
60.00000000000,0.0000
61.00000000000,0.0000
62.00000000000,0.0000
63.00000000000,0.0000
64.00000000000,0.0000
65.00000000000,0.0000
66.00000000000,0.0000
67.00000000000,0.0000
68.00000000000,0.0000
69.00000000000,778.43
70.00000000000,0.0000
71.00000000000,0.0000
72.00000000000,0.0000
73.00000000000,0.0000
74.00000000000,0.0000
75.00000000000,0.0000
76.00000000000,0.0000
77.00000000000,0.0000
78.00000000000,0.0000
79.00000000000,0.0000
80.00000000000,0.0000
81.00000000000,0.0000
82.00000000000,446.67
83.00000000000,0.0000
84.00000000000,0.0000
85.00000000000,0.0000
86.00000000000,0.0000
87.00000000000,0.0000
88.00000000000,0.0000
89.00000000000,0.0000
90.00000000000,0.0000
91.00000000000,2.8531
92.00000000000,6.9710
93.00000000000,1938.4
94.00000000000,30.640
95.00000000000,0.0000
96.00000000000,0.0000
97.00000000000,0.0000
98.00000000000,0.0000
99.00000000000,0.0000
100.0000000000,0.0000
101.0000000000,0.0000
102.0000000000,0.0000
103.0000000000,0.0000
104.0000000000,0.0000
105.0000000000,0.0000
106.0000000000,0.0000
107.0000000000,0.0000
108.0000000000,1117.7
109.0000000000,0.0000
110.0000000000,0.0000
111.0000000000,0.0000
112.0000000000,0.0000
113.0000000000,0.0000
114.0000000000,0.0000
115.0000000000,0.0000
116.0000000000,0.0000
117.0000000000,0.0000
118.0000000000,3675.8
119.0000000000,6271.9
120.0000000000,0.0000
121.0000000000,0.0000
122.0000000000,2359.3
123.0000000000,0.0000
124.0000000000,0.0000
125.0000000000,0.0000
126.0000000000,0.0000
127.0000000000,0.0000
128.0000000000,0.0000
129.0000000000,0.0000
130.0000000000,1193.1
131.0000000000,1472.4
132.0000000000,0.0000
133.0000000000,0.0000
134.0000000000,0.0000
135.0000000000,1943.6
136.0000000000,0.0000
137.0000000000,0.0000
138.0000000000,0.0000
139.0000000000,0.0000
140.0000000000,0.0000
141.0000000000,0.0000
142.0000000000,0.0000
143.0000000000,0.0000
144.0000000000,4386.2
145.0000000000,360.16
146.0000000000,6845.6
147.0000000000,0.0000
148.0000000000,0.0000
149.0000000000,956.26
150.0000000000,7.4573
151.0000000000,0.0000
152.0000000000,0.0000
153.0000000000,0.0000
154.0000000000,143.26
155.0000000000,0.0000
156.0000000000,0.0000
157.0000000000,0.0000
158.0000000000,36.768
159.0000000000,1546.7
160.0000000000,0.0000
161.0000000000,5.2196
162.0000000000,0.0000
163.0000000000,0.0000
164.0000000000,0.0000
165.0000000000,983.44
166.0000000000,8786.2
167.0000000000,655.44
168.0000000000,0.0000
169.0000000000,652.77
170.0000000000,192.21
171.0000000000,0.0000
172.0000000000,0.0000
173.0000000000,0.0000
174.0000000000,0.0000
175.0000000000,0.0000
176.0000000000,0.0000
177.0000000000,0.0000
178.0000000000,0.0000
179.0000000000,0.0000
180.0000000000,0.0000
181.0000000000,2178.9
182.0000000000,23.143
183.0000000000,488.36
184.0000000000,0.0000
185.0000000000,0.0000
186.0000000000,0.0000
187.0000000000,0.0000
188.0000000000,0.0000
189.0000000000,0.0000
190.0000000000,0.0000
191.0000000000,0.0000
192.0000000000,0.0000
193.0000000000,0.0000
194.0000000000,0.0000
195.0000000000,0.0000
196.0000000000,551.97
197.0000000000,5728.2
198.0000000000,3023.5
199.0000000000,563.91
200.0000000000,915.04
201.0000000000,13.913
202.0000000000,152.40
203.0000000000,241.77
204.0000000000,0.0000
205.0000000000,0.0000
206.0000000000,0.0000
207.0000000000,0.0000
208.0000000000,253.98
209.0000000000,0.0000
210.0000000000,848.57
211.0000000000,0.0000
212.0000000000,0.0000
213.0000000000,0.0000
214.0000000000,12.624
215.0000000000,0.0000
216.0000000000,0.0000
217.0000000000,0.0000
218.0000000000,0.0000
219.0000000000,0.0000
220.0000000000,0.0000
221.0000000000,0.0000
222.0000000000,0.0000
223.0000000000,50.368
224.0000000000,276.42
225.0000000000,0.0000
226.0000000000,0.0000
227.0000000000,0.0000
228.0000000000,2.6547
229.0000000000,0.33931E-01
230.0000000000,0.0000
231.0000000000,4.1530
232.0000000000,0.0000
233.0000000000,0.0000
234.0000000000,172.84
235.0000000000,0.0000
236.0000000000,4583.1
237.0000000000,102.86
238.0000000000,662.05
239.0000000000,5919.0
240.0000000000,4811.3
241.0000000000,0.0000
242.0000000000,0.0000
243.0000000000,0.0000
244.0000000000,0.0000
245.0000000000,2.4855
246.0000000000,2079.0
247.0000000000,0.0000
248.0000000000,1624.9
249.0000000000,988.63
250.0000000000,0.0000
251.0000000000,0.0000
252.0000000000,1317.6
253.0000000000,221.33
254.0000000000,653.66
255.0000000000,6.4219
256.0000000000,0.0000
257.0000000000,0.0000
258.0000000000,0.0000
259.0000000000,0.0000
260.0000000000,1118.0
261.0000000000,2184.5
262.0000000000,511.81
263.0000000000,13083.
264.0000000000,10638.
265.0000000000,0.0000
266.0000000000,0.0000
267.0000000000,0.0000
268.0000000000,0.0000
269.0000000000,0.0000
270.0000000000,0.0000
271.0000000000,0.0000
272.0000000000,1777.3
273.0000000000,0.0000
274.0000000000,0.0000
275.0000000000,0.0000
276.0000000000,0.0000
277.0000000000,0.0000
278.0000000000,0.0000
279.0000000000,17.697
280.0000000000,0.0000
281.0000000000,0.0000
282.0000000000,0.0000
283.0000000000,0.0000
284.0000000000,0.0000
285.0000000000,0.0000
286.0000000000,47.572
287.0000000000,1592.0
288.0000000000,2899.5
289.0000000000,8821.5
290.0000000000,217.33
291.0000000000,0.0000
292.0000000000,41.666
293.0000000000,0.0000
294.0000000000,0.0000
295.0000000000,0.0000
296.0000000000,0.0000
297.0000000000,0.0000
298.0000000000,0.0000
299.0000000000,0.0000
300.0000000000,0.0000
301.0000000000,0.0000
302.0000000000,0.0000
303.0000000000,0.0000
304.0000000000,73.397
305.0000000000,0.0000
306.0000000000,0.0000
307.0000000000,0.0000
308.0000000000,1139.6
309.0000000000,317.40
310.0000000000,957.80
311.0000000000,789.81
312.0000000000,0.0000
313.0000000000,920.31
314.0000000000,0.0000
315.0000000000,0.0000
316.0000000000,189.01
317.0000000000,45.836
318.0000000000,0.0000
319.0000000000,0.0000
320.0000000000,0.0000
321.0000000000,0.0000
322.0000000000,0.0000
323.0000000000,0.0000
324.0000000000,0.0000
325.0000000000,0.0000
326.0000000000,361.66
327.0000000000,348.75
328.0000000000,2349.3
329.0000000000,1884.8
330.0000000000,40.930
331.0000000000,0.0000
332.0000000000,0.0000
333.0000000000,0.0000
334.0000000000,0.0000
335.0000000000,0.0000
336.0000000000,0.0000
337.0000000000,0.0000
338.0000000000,0.0000
339.0000000000,0.0000
340.0000000000,449.24
341.0000000000,1.6340
342.0000000000,0.0000
343.0000000000,0.0000
344.0000000000,0.0000
345.0000000000,0.0000
346.0000000000,0.0000
347.0000000000,0.0000
348.0000000000,0.0000
349.0000000000,0.0000
350.0000000000,0.0000
351.0000000000,0.0000
352.0000000000,0.0000
353.0000000000,0.0000
354.0000000000,0.0000
355.0000000000,1733.9
356.0000000000,652.84
357.0000000000,0.0000
358.0000000000,0.0000
359.0000000000,0.0000
360.0000000000,574.98
361.0000000000,1162.8
362.0000000000,1010.6
363.0000000000,0.0000
364.0000000000,0.0000
365.0000000000,0.0000
366.0000000000,0.0000
367.0000000000,0.0000
368.0000000000,0.0000
369.0000000000,0.0000
370.0000000000,0.0000
371.0000000000,0.0000
372.0000000000,0.0000
373.0000000000,0.0000
374.0000000000,0.0000
375.0000000000,0.0000
376.0000000000,0.0000
377.0000000000,0.0000
378.0000000000,0.0000
379.0000000000,0.0000
380.0000000000,0.0000
381.0000000000,0.0000
382.0000000000,0.0000
383.0000000000,0.0000
384.0000000000,0.0000
385.0000000000,0.0000
386.0000000000,0.0000
387.0000000000,0.0000
388.0000000000,0.0000
389.0000000000,149.95
390.0000000000,0.0000
391.0000000000,0.0000
392.0000000000,0.0000
393.0000000000,0.0000
394.0000000000,0.0000
395.0000000000,0.0000
396.0000000000,0.0000
397.0000000000,0.0000
398.0000000000,0.0000
399.0000000000,5.1474
400.0000000000,0.0000
401.0000000000,0.0000
402.0000000000,0.0000
403.0000000000,0.0000
404.0000000000,0.0000
405.0000000000,0.0000
406.0000000000,0.0000
407.0000000000,0.0000
408.0000000000,0.0000
409.0000000000,0.0000
410.0000000000,0.0000
411.0000000000,0.0000
412.0000000000,0.0000
413.0000000000,0.0000
414.0000000000,0.0000
415.0000000000,0.0000
416.0000000000,0.0000
417.0000000000,0.0000
418.0000000000,0.0000
419.0000000000,0.0000
420.0000000000,0.0000
421.0000000000,102.71
422.0000000000,1505.8
423.0000000000,461.07
424.0000000000,0.0000
425.0000000000,0.0000
426.0000000000,42.453
427.0000000000,0.0000
428.0000000000,4.3267
429.0000000000,0.0000
430.0000000000,0.0000
431.0000000000,0.0000
432.0000000000,0.0000
433.0000000000,0.0000
434.0000000000,63.381
435.0000000000,0.13997
436.0000000000,0.0000
437.0000000000,0.0000
438.0000000000,0.0000
439.0000000000,0.0000
440.0000000000,0.0000
441.0000000000,0.0000
442.0000000000,0.0000
443.0000000000,0.0000
444.0000000000,0.0000
445.0000000000,0.0000
446.0000000000,0.0000
447.0000000000,0.0000
448.0000000000,337.78
449.0000000000,0.0000
450.0000000000,0.0000
451.0000000000,57.941
452.0000000000,0.0000
453.0000000000,0.0000
454.0000000000,0.0000
455.0000000000,0.0000
456.0000000000,0.0000
457.0000000000,0.0000
458.0000000000,0.0000
459.0000000000,1270.7
460.0000000000,0.0000
461.0000000000,57.868
462.0000000000,9.6503
463.0000000000,140.84
464.0000000000,0.0000
465.0000000000,0.0000
466.0000000000,0.0000
467.0000000000,0.0000
468.0000000000,0.0000
469.0000000000,18.536
470.0000000000,0.0000
471.0000000000,0.0000
472.0000000000,0.0000
473.0000000000,0.0000
474.0000000000,0.0000
475.0000000000,161.30
476.0000000000,0.0000
477.0000000000,0.21905
478.0000000000,0.0000
479.0000000000,0.0000
480.0000000000,0.0000
481.0000000000,0.0000
482.0000000000,0.0000
483.0000000000,0.0000
484.0000000000,0.0000
485.0000000000,0.0000
486.0000000000,0.0000
487.0000000000,0.0000
488.0000000000,0.0000
489.0000000000,0.0000
490.0000000000,0.0000
491.0000000000,0.0000
492.0000000000,967.81
493.0000000000,0.25710E-01
494.0000000000,444.80
495.0000000000,851.58
496.0000000000,0.0000
497.0000000000,38.244
498.0000000000,936.06
499.0000000000,214.89
500.0000000000,0.0000
501.0000000000,0.0000
502.0000000000,0.0000
503.0000000000,0.0000
504.0000000000,0.0000
505.0000000000,0.0000
506.0000000000,0.0000
507.0000000000,0.0000
508.0000000000,369.59
509.0000000000,15.624
510.0000000000,919.06
511.0000000000,6137.9
512.0000000000,392.76
513.0000000000,0.0000
514.0000000000,0.0000
515.0000000000,0.0000
516.0000000000,0.0000
517.0000000000,0.0000
518.0000000000,0.0000
519.0000000000,0.0000
520.0000000000,0.0000
521.0000000000,0.0000
522.0000000000,0.0000
523.0000000000,0.0000
524.0000000000,0.0000
525.0000000000,90.078
526.0000000000,64.470
527.0000000000,0.0000
528.0000000000,196.03
529.0000000000,1246.0
530.0000000000,2318.4
531.0000000000,26.375
532.0000000000,0.0000
533.0000000000,0.0000
534.0000000000,0.0000
535.0000000000,0.10957
536.0000000000,13476.
537.0000000000,5684.7
538.0000000000,1890.8
539.0000000000,0.0000
540.0000000000,108.66
541.0000000000,4909.3
542.0000000000,0.0000
543.0000000000,0.0000
544.0000000000,66.650
545.0000000000,0.0000
546.0000000000,0.0000
547.0000000000,0.0000
548.0000000000,0.0000
549.0000000000,12.747
550.0000000000,0.0000
551.0000000000,0.0000
552.0000000000,0.0000
553.0000000000,0.0000
554.0000000000,0.0000
555.0000000000,0.0000
556.0000000000,59.792
557.0000000000,73.526
558.0000000000,1020.7
559.0000000000,0.0000
560.0000000000,0.0000
561.0000000000,0.0000
562.0000000000,1338.5
563.0000000000,1607.4
564.0000000000,1193.1
565.0000000000,0.0000
566.0000000000,0.0000
567.0000000000,0.0000
568.0000000000,0.0000
569.0000000000,0.0000
570.0000000000,0.0000
571.0000000000,568.43
572.0000000000,0.0000
573.0000000000,0.0000
574.0000000000,0.0000
575.0000000000,0.0000
576.0000000000,0.0000
577.0000000000,0.0000
578.0000000000,3.1775
579.0000000000,2389.8
580.0000000000,6246.7
581.0000000000,0.0000
582.0000000000,0.0000
583.0000000000,0.0000
584.0000000000,0.0000
585.0000000000,0.0000
586.0000000000,0.0000
587.0000000000,0.0000
588.0000000000,0.0000
589.0000000000,643.52
590.0000000000,1510.8
591.0000000000,0.0000
592.0000000000,0.0000
593.0000000000,0.72141E-01
594.0000000000,379.72
595.0000000000,1908.7
596.0000000000,2362.4
597.0000000000,8.6521
598.0000000000,0.0000
599.0000000000,0.0000
600.0000000000,0.0000
601.0000000000,0.0000
602.0000000000,0.0000
603.0000000000,0.0000
604.0000000000,0.10480
605.0000000000,49.351
606.0000000000,0.0000
607.0000000000,288.83
608.0000000000,77.441
609.0000000000,0.0000
610.0000000000,0.0000
611.0000000000,0.0000
612.0000000000,35.552
613.0000000000,1901.2
614.0000000000,535.35
615.0000000000,10.064
616.0000000000,1413.2
617.0000000000,5.1823
618.0000000000,0.0000
619.0000000000,0.0000
620.0000000000,47.542
621.0000000000,551.19
622.0000000000,434.30
623.0000000000,40.440
624.0000000000,0.0000
625.0000000000,323.41
626.0000000000,8.0902
627.0000000000,3324.0
628.0000000000,290.62
629.0000000000,1628.6
630.0000000000,967.30
631.0000000000,0.0000
632.0000000000,0.0000
633.0000000000,33.627
634.0000000000,84.070
635.0000000000,7252.3
636.0000000000,1275.7
637.0000000000,0.0000
638.0000000000,0.0000
639.0000000000,0.0000
640.0000000000,0.0000
641.0000000000,0.0000
642.0000000000,0.0000
643.0000000000,0.0000
644.0000000000,0.0000
645.0000000000,0.0000
646.0000000000,0.0000
647.0000000000,0.0000
648.0000000000,0.0000
649.0000000000,3006.3
650.0000000000,0.0000
651.0000000000,0.0000
652.0000000000,0.0000
653.0000000000,0.0000
654.0000000000,0.0000
655.0000000000,0.0000
656.0000000000,0.0000
657.0000000000,0.0000
658.0000000000,0.22293
659.0000000000,124.37
660.0000000000,567.99
661.0000000000,1707.5
662.0000000000,0.0000
663.0000000000,0.0000
664.0000000000,0.0000
665.0000000000,0.0000
666.0000000000,0.0000
667.0000000000,0.0000
668.0000000000,0.26199E-01
669.0000000000,0.26199E-01
670.0000000000,0.0000
671.0000000000,0.0000
672.0000000000,0.0000
673.0000000000,0.0000
674.0000000000,10103.
675.0000000000,5596.0
676.0000000000,188.65
677.0000000000,127.34
678.0000000000,0.0000
679.0000000000,0.0000
680.0000000000,0.0000
681.0000000000,0.0000
682.0000000000,0.0000
683.0000000000,0.0000
684.0000000000,0.0000
685.0000000000,0.0000
686.0000000000,0.0000
687.0000000000,0.0000
688.0000000000,0.0000
689.0000000000,0.0000
690.0000000000,0.0000
691.0000000000,1.4237
692.0000000000,909.50
693.0000000000,0.0000
694.0000000000,0.0000
695.0000000000,0.0000
696.0000000000,0.0000
697.0000000000,0.0000
698.0000000000,0.0000
699.0000000000,0.0000
700.0000000000,0.0000
701.0000000000,0.0000
702.0000000000,0.0000
703.0000000000,0.0000
704.0000000000,0.0000
705.0000000000,0.0000
706.0000000000,0.0000
707.0000000000,0.0000
708.0000000000,0.0000
709.0000000000,12.352
710.0000000000,53.007
711.0000000000,0.0000
712.0000000000,0.0000
713.0000000000,0.0000
714.0000000000,0.0000
715.0000000000,0.0000
716.0000000000,0.0000
717.0000000000,0.0000
718.0000000000,102.97
719.0000000000,0.0000
720.0000000000,0.0000
721.0000000000,0.0000
722.0000000000,97.909
723.0000000000,123.56
724.0000000000,0.0000
725.0000000000,0.0000
726.0000000000,0.0000
727.0000000000,3901.3
728.0000000000,174.27
729.0000000000,0.0000
730.0000000000,224.54
731.0000000000,740.36
732.0000000000,1182.8
733.0000000000,1338.7
734.0000000000,0.0000
735.0000000000,0.0000
736.0000000000,0.0000
737.0000000000,0.0000
738.0000000000,0.0000
739.0000000000,88.290
740.0000000000,1882.8
741.0000000000,192.75
742.0000000000,6.9230
743.0000000000,0.0000
744.0000000000,0.0000
745.0000000000,0.0000
746.0000000000,0.0000
747.0000000000,0.0000
748.0000000000,0.0000
749.0000000000,0.0000
750.0000000000,0.0000
751.0000000000,0.0000
752.0000000000,1248.7
753.0000000000,1439.5
754.0000000000,91.004
755.0000000000,0.0000
756.0000000000,0.0000
757.0000000000,0.0000
758.0000000000,0.0000
759.0000000000,0.0000
760.0000000000,0.0000
761.0000000000,1137.7
762.0000000000,1574.5
763.0000000000,0.0000
764.0000000000,0.0000
765.0000000000,77.651
766.0000000000,0.0000
767.0000000000,0.0000
768.0000000000,0.0000
769.0000000000,0.0000
770.0000000000,0.0000
771.0000000000,0.0000
772.0000000000,0.0000
773.0000000000,0.0000
774.0000000000,0.0000
775.0000000000,0.0000
776.0000000000,0.0000
777.0000000000,25.216
778.0000000000,126.34
779.0000000000,0.0000
780.0000000000,0.0000
781.0000000000,0.0000
782.0000000000,0.0000
783.0000000000,0.0000
784.0000000000,0.0000
785.0000000000,0.0000
786.0000000000,0.0000
787.0000000000,0.0000
788.0000000000,0.0000
789.0000000000,469.58
790.0000000000,133.66
791.0000000000,55.495
792.0000000000,0.0000
793.0000000000,0.0000
794.0000000000,1725.3
795.0000000000,0.0000
796.0000000000,0.0000
797.0000000000,563.61
798.0000000000,128.91
799.0000000000,226.31
800.0000000000,0.0000
801.0000000000,0.0000
802.0000000000,0.0000
803.0000000000,0.0000
804.0000000000,0.0000
805.0000000000,0.0000
806.0000000000,0.0000
807.0000000000,369.99
808.0000000000,37.500
809.0000000000,1934.8
810.0000000000,7024.1
811.0000000000,4016.7
812.0000000000,0.0000
813.0000000000,0.0000
814.0000000000,0.0000
815.0000000000,242.78
816.0000000000,0.0000
817.0000000000,0.0000
818.0000000000,0.0000
819.0000000000,0.0000
820.0000000000,0.0000
821.0000000000,0.0000
822.0000000000,0.0000
823.0000000000,0.0000
824.0000000000,0.0000
825.0000000000,0.0000
826.0000000000,347.81
827.0000000000,0.0000
828.0000000000,93.371
829.0000000000,822.93
830.0000000000,3.0689
831.0000000000,0.0000
832.0000000000,564.28
833.0000000000,3080.8
834.0000000000,0.0000
835.0000000000,0.0000
836.0000000000,1600.2
837.0000000000,386.95
838.0000000000,2390.3
839.0000000000,61.491
840.0000000000,0.0000
841.0000000000,0.0000
842.0000000000,0.0000
843.0000000000,0.0000
844.0000000000,1745.0
845.0000000000,0.0000
846.0000000000,0.0000
847.0000000000,2930.3
848.0000000000,0.0000
849.0000000000,0.0000
850.0000000000,0.0000
851.0000000000,0.0000
852.0000000000,0.0000
853.0000000000,0.0000
854.0000000000,0.0000
855.0000000000,24.723
856.0000000000,0.0000
857.0000000000,68.672
858.0000000000,0.0000
859.0000000000,0.0000
860.0000000000,0.66706E-01
861.0000000000,9096.2
862.0000000000,6700.5
863.0000000000,4921.4
864.0000000000,1873.2
865.0000000000,999.26
866.0000000000,3778.2
867.0000000000,6738.6
868.0000000000,0.0000
869.0000000000,34.838
870.0000000000,0.0000
871.0000000000,2952.7
872.0000000000,610.84
873.0000000000,160.43
874.0000000000,1748.1
875.0000000000,161.25
876.0000000000,734.86
877.0000000000,0.0000
878.0000000000,0.0000
879.0000000000,7620.3
880.0000000000,132.84
881.0000000000,5926.2
882.0000000000,0.0000
883.0000000000,0.0000
884.0000000000,0.0000
885.0000000000,0.0000
886.0000000000,0.0000
887.0000000000,0.0000
888.0000000000,0.0000
889.0000000000,0.0000
890.0000000000,0.0000
891.0000000000,0.0000
892.0000000000,0.0000
893.0000000000,0.0000
894.0000000000,620.80
895.0000000000,5023.6
896.0000000000,555.69
897.0000000000,2391.9
898.0000000000,1006.9
899.0000000000,139.75
900.0000000000,54.751
901.0000000000,2329.2
902.0000000000,246.83
903.0000000000,0.0000
904.0000000000,586.45
905.0000000000,30.026
906.0000000000,0.0000
907.0000000000,0.0000
908.0000000000,2991.8
909.0000000000,2715.4
910.0000000000,145.42
911.0000000000,12.643
912.0000000000,705.73
913.0000000000,0.0000
914.0000000000,0.0000
915.0000000000,0.0000
916.0000000000,0.0000
917.0000000000,0.0000
918.0000000000,20.421
919.0000000000,3058.3
920.0000000000,0.0000
921.0000000000,0.0000
922.0000000000,0.0000
923.0000000000,0.0000
924.0000000000,0.0000
925.0000000000,0.0000
926.0000000000,0.0000
927.0000000000,0.0000
928.0000000000,0.0000
929.0000000000,0.0000
930.0000000000,0.0000
931.0000000000,0.0000
932.0000000000,0.0000
933.0000000000,0.0000
934.0000000000,0.0000
935.0000000000,0.0000
936.0000000000,0.0000
937.0000000000,0.0000
938.0000000000,0.0000
939.0000000000,0.0000
940.0000000000,0.0000
941.0000000000,0.0000
942.0000000000,0.0000
943.0000000000,847.35
944.0000000000,860.61
945.0000000000,0.0000
946.0000000000,0.0000
947.0000000000,0.0000
948.0000000000,0.0000
949.0000000000,0.0000
950.0000000000,0.0000
951.0000000000,0.0000
952.0000000000,0.0000
953.0000000000,0.0000
954.0000000000,0.0000
955.0000000000,854.17
956.0000000000,642.45
957.0000000000,1295.4
958.0000000000,1866.6
959.0000000000,0.0000
960.0000000000,0.0000
961.0000000000,0.0000
962.0000000000,2583.2
963.0000000000,1133.3
964.0000000000,0.0000
965.0000000000,0.0000
966.0000000000,0.0000
967.0000000000,0.0000
968.0000000000,493.00
969.0000000000,620.95
970.0000000000,0.0000
971.0000000000,0.0000
972.0000000000,0.0000
973.0000000000,334.94
974.0000000000,0.0000
975.0000000000,0.0000
976.0000000000,0.0000
977.0000000000,0.0000
978.0000000000,0.0000
979.0000000000,0.0000
980.0000000000,0.0000
981.0000000000,0.0000
982.0000000000,0.0000
983.0000000000,1497.9
984.0000000000,5.8475
985.0000000000,877.21
986.0000000000,0.0000
987.0000000000,0.0000
988.0000000000,0.0000
989.0000000000,0.0000
990.0000000000,0.0000
991.0000000000,0.0000
992.0000000000,0.0000
993.0000000000,0.0000
994.0000000000,0.0000
995.0000000000,0.0000
996.0000000000,0.0000
997.0000000000,0.0000
998.0000000000,0.0000
999.0000000000,0.0000
1000.000000000,614.88
1001.000000000,0.0000
1002.000000000,0.0000
1003.000000000,0.0000
1004.000000000,0.0000
1005.000000000,0.0000
1006.000000000,0.0000
1007.000000000,0.0000
1008.000000000,0.0000
1009.000000000,17.919
1010.000000000,0.0000
1011.000000000,0.0000
1012.000000000,7036.3
1013.000000000,1098.0
1014.000000000,0.0000
1015.000000000,0.0000
1016.000000000,0.0000
1017.000000000,0.0000
1018.000000000,0.0000
1019.000000000,0.0000
1020.000000000,0.0000
1021.000000000,0.0000
1022.000000000,0.0000
1023.000000000,0.0000
1024.000000000,0.0000
1025.000000000,435.41
1026.000000000,770.69
1027.000000000,14579.
1028.000000000,6396.0
1029.000000000,0.0000
1030.000000000,0.0000
1031.000000000,0.0000
1032.000000000,0.0000
1033.000000000,569.92
1034.000000000,8508.7
1035.000000000,0.0000
1036.000000000,0.0000
1037.000000000,0.0000
1038.000000000,0.0000
1039.000000000,0.0000
1040.000000000,0.0000
1041.000000000,358.09
1042.000000000,323.53
1043.000000000,0.0000
1044.000000000,0.0000
1045.000000000,0.0000
1046.000000000,0.0000
1047.000000000,0.0000
1048.000000000,176.78
1049.000000000,615.14
1050.000000000,111.47
1051.000000000,202.98
1052.000000000,0.0000
1053.000000000,0.0000
1054.000000000,0.0000
1055.000000000,0.0000
1056.000000000,0.0000
1057.000000000,0.0000
1058.000000000,0.0000
1059.000000000,0.0000
1060.000000000,263.23
1061.000000000,1257.1
1062.000000000,5288.2
1063.000000000,227.35
1064.000000000,1.0046
1065.000000000,0.0000
1066.000000000,0.0000
1067.000000000,0.0000
1068.000000000,0.0000
1069.000000000,0.0000
1070.000000000,0.0000
1071.000000000,0.0000
1072.000000000,0.0000
1073.000000000,0.0000
1074.000000000,0.0000
1075.000000000,0.0000
1076.000000000,0.0000
1077.000000000,6203.6
1078.000000000,0.0000
1079.000000000,0.0000
1080.000000000,0.0000
1081.000000000,0.0000
1082.000000000,0.0000
1083.000000000,0.0000
1084.000000000,0.79079
1085.000000000,0.21913
1086.000000000,0.0000
1087.000000000,0.0000
1088.000000000,0.0000
1089.000000000,0.0000
1090.000000000,0.0000
1091.000000000,5257.9
1092.000000000,1078.3
1093.000000000,0.0000
1094.000000000,0.0000
1095.000000000,0.0000
1096.000000000,0.0000
1097.000000000,68.462
1098.000000000,955.95
1099.000000000,0.0000
1100.000000000,0.0000
1101.000000000,0.0000
1102.000000000,0.0000
1103.000000000,0.0000
1104.000000000,0.0000
1105.000000000,0.0000
1106.000000000,0.0000
1107.000000000,0.0000
1108.000000000,0.0000
1109.000000000,0.0000
1110.000000000,0.0000
1111.000000000,0.0000
1112.000000000,0.0000
1113.000000000,0.0000
1114.000000000,0.0000
1115.000000000,0.0000
1116.000000000,0.0000
1117.000000000,0.0000
1118.000000000,0.0000
1119.000000000,0.0000
1120.000000000,0.0000
1121.000000000,0.0000
1122.000000000,3207.1
1123.000000000,0.0000
1124.000000000,0.0000
1125.000000000,0.0000
1126.000000000,0.0000
1127.000000000,0.0000
1128.000000000,0.0000
1129.000000000,0.0000
1130.000000000,0.0000
1131.000000000,0.0000
1132.000000000,0.0000
1133.000000000,0.0000
1134.000000000,0.0000
1135.000000000,0.0000
1136.000000000,0.0000
1137.000000000,0.0000
1138.000000000,0.0000
1139.000000000,0.0000
1140.000000000,0.0000
1141.000000000,0.0000
1142.000000000,0.0000
1143.000000000,0.0000
1144.000000000,0.0000
1145.000000000,0.0000
1146.000000000,0.0000
1147.000000000,0.0000
1148.000000000,1224.5
1149.000000000,3390.3
1150.000000000,0.0000
1151.000000000,0.0000
1152.000000000,0.0000
1153.000000000,0.0000
1154.000000000,0.0000
1155.000000000,0.0000
1156.000000000,0.0000
1157.000000000,0.0000
1158.000000000,0.0000
1159.000000000,0.0000
1160.000000000,0.0000
1161.000000000,0.0000
1162.000000000,0.0000
1163.000000000,5655.4
1164.000000000,3589.6
1165.000000000,5355.6
1166.000000000,5312.6
1167.000000000,3249.3
1168.000000000,0.0000
1169.000000000,0.0000
1170.000000000,0.0000
1171.000000000,0.0000
1172.000000000,97.242
1173.000000000,0.0000
1174.000000000,2613.3
1175.000000000,0.0000
1176.000000000,0.0000
1177.000000000,0.0000
1178.000000000,0.0000
1179.000000000,346.12
1180.000000000,0.0000
1181.000000000,0.0000
1182.000000000,0.0000
1183.000000000,0.0000
1184.000000000,0.0000
1185.000000000,0.0000
1186.000000000,0.0000
1187.000000000,56.063
1188.000000000,0.0000
1189.000000000,0.0000
1190.000000000,0.0000
1191.000000000,0.0000
1192.000000000,0.0000
1193.000000000,0.0000
1194.000000000,0.0000
1195.000000000,0.0000
1196.000000000,0.0000
1197.000000000,89.671
1198.000000000,0.0000
1199.000000000,2336.7
1200.000000000,0.0000
1201.000000000,0.0000
1202.000000000,0.0000
1203.000000000,15507.
1204.000000000,3409.9
1205.000000000,87.464
1206.000000000,83.633
1207.000000000,20.529
1208.000000000,53.659
1209.000000000,0.0000
1210.000000000,243.39
1211.000000000,0.0000
1212.000000000,0.0000
1213.000000000,1534.6
1214.000000000,0.0000
1215.000000000,0.0000
1216.000000000,45.429
1217.000000000,0.0000
1218.000000000,58.498
1219.000000000,0.0000
1220.000000000,0.0000
1221.000000000,0.0000
1222.000000000,0.0000
1223.000000000,0.0000
1224.000000000,0.0000
1225.000000000,501.56
1226.000000000,0.0000
1227.000000000,0.0000
1228.000000000,0.0000
1229.000000000,64.334
1230.000000000,5.8804
1231.000000000,802.99
1232.000000000,501.81
1233.000000000,14.806
1234.000000000,1877.2
1235.000000000,4910.2
1236.000000000,982.53
1237.000000000,0.0000
1238.000000000,0.0000
1239.000000000,0.0000
1240.000000000,0.21275
1241.000000000,0.0000
1242.000000000,0.0000
1243.000000000,42.726
1244.000000000,0.0000
1245.000000000,0.35495
1246.000000000,220.55
1247.000000000,0.0000
1248.000000000,560.42
1249.000000000,10071.
1250.000000000,2210.2
1251.000000000,203.60
1252.000000000,0.85702E-01
1253.000000000,0.0000
1254.000000000,0.0000
1255.000000000,0.0000
1256.000000000,0.0000
1257.000000000,0.0000
1258.000000000,0.0000
1259.000000000,0.0000
1260.000000000,105.28
1261.000000000,0.0000
1262.000000000,0.0000
1263.000000000,0.0000
1264.000000000,0.0000
1265.000000000,0.0000
1266.000000000,0.0000
1267.000000000,2227.3
1268.000000000,0.0000
1269.000000000,0.0000
1270.000000000,0.0000
1271.000000000,0.0000
1272.000000000,0.0000
1273.000000000,2148.2
1274.000000000,16846.
1275.000000000,595.53
1276.000000000,189.19
1277.000000000,0.0000
1278.000000000,13.478
1279.000000000,0.0000
1280.000000000,0.0000
1281.000000000,0.0000
1282.000000000,0.0000
1283.000000000,0.0000
1284.000000000,0.0000
1285.000000000,0.0000
1286.000000000,0.0000
1287.000000000,19.659
1288.000000000,0.0000
1289.000000000,0.0000
1290.000000000,0.0000
1291.000000000,0.0000
1292.000000000,0.0000
1293.000000000,0.0000
1294.000000000,0.0000
1295.000000000,0.0000
1296.000000000,0.0000
1297.000000000,0.0000
1298.000000000,0.0000
1299.000000000,0.0000
1300.000000000,0.0000
1301.000000000,0.0000
1302.000000000,0.0000
1303.000000000,55.886
1304.000000000,1753.3
1305.000000000,161.98
1306.000000000,0.95602
1307.000000000,73.160
1308.000000000,0.0000
1309.000000000,0.0000
1310.000000000,0.0000
1311.000000000,0.0000
1312.000000000,0.0000
1313.000000000,0.0000
1314.000000000,0.0000
1315.000000000,0.0000
1316.000000000,0.0000
1317.000000000,0.0000
1318.000000000,0.0000
1319.000000000,0.0000
1320.000000000,0.0000
1321.000000000,6179.1
1322.000000000,5344.4
1323.000000000,2039.1
1324.000000000,410.38
1325.000000000,3765.4
1326.000000000,1161.5
1327.000000000,448.32
1328.000000000,12990.
1329.000000000,1634.5
1330.000000000,2510.0
1331.000000000,3075.1
1332.000000000,0.0000
1333.000000000,406.32
1334.000000000,0.0000
1335.000000000,1.5004
1336.000000000,211.13
1337.000000000,938.03
1338.000000000,417.15
1339.000000000,880.85
1340.000000000,520.55
1341.000000000,520.63
1342.000000000,1867.9
1343.000000000,31.089
1344.000000000,0.0000
1345.000000000,14.792
1346.000000000,0.0000
1347.000000000,0.0000
1348.000000000,0.0000
1349.000000000,0.0000
1350.000000000,656.10
1351.000000000,0.0000
1352.000000000,1696.6
1353.000000000,157.49
1354.000000000,753.31
1355.000000000,0.0000
1356.000000000,0.0000
1357.000000000,0.0000
1358.000000000,0.0000
1359.000000000,0.0000
1360.000000000,0.0000
1361.000000000,0.0000
1362.000000000,0.0000
1363.000000000,0.0000
1364.000000000,8153.6
1365.000000000,18740.
1366.000000000,2053.6
1367.000000000,0.0000
1368.000000000,0.0000
1369.000000000,0.0000
1370.000000000,0.0000
1371.000000000,0.36500
1372.000000000,0.0000
1373.000000000,0.0000
1374.000000000,0.0000
1375.000000000,0.0000
1376.000000000,0.0000
1377.000000000,40.927
1378.000000000,0.0000
1379.000000000,0.0000
1380.000000000,0.0000
1381.000000000,0.0000
1382.000000000,0.0000
1383.000000000,0.0000
1384.000000000,0.0000
1385.000000000,0.0000
1386.000000000,0.0000
1387.000000000,0.0000
1388.000000000,0.0000
1389.000000000,0.0000
1390.000000000,34.493
1391.000000000,0.0000
1392.000000000,0.0000
1393.000000000,0.0000
1394.000000000,0.0000
1395.000000000,0.0000
1396.000000000,0.0000
1397.000000000,0.0000
1398.000000000,0.0000
1399.000000000,0.0000
1400.000000000,0.0000
1401.000000000,0.0000
1402.000000000,0.0000
1403.000000000,0.0000
1404.000000000,3576.6
1405.000000000,127.54
1406.000000000,60.647
1407.000000000,478.68
1408.000000000,0.0000
1409.000000000,0.0000
1410.000000000,5372.1
1411.000000000,165.32
1412.000000000,0.0000
1413.000000000,0.0000
1414.000000000,0.0000
1415.000000000,0.0000
1416.000000000,0.0000
1417.000000000,0.0000
1418.000000000,0.0000
1419.000000000,0.0000
1420.000000000,0.0000
1421.000000000,0.0000
1422.000000000,0.0000
1423.000000000,0.0000
1424.000000000,0.0000
1425.000000000,0.0000
1426.000000000,486.23
1427.000000000,0.0000
1428.000000000,0.0000
1429.000000000,0.0000
1430.000000000,0.0000
1431.000000000,0.0000
1432.000000000,0.0000
1433.000000000,2053.5
1434.000000000,3479.4
1435.000000000,11700.
1436.000000000,1148.7
1437.000000000,0.0000
1438.000000000,0.0000
1439.000000000,0.0000
1440.000000000,0.0000
1441.000000000,0.0000
1442.000000000,0.0000
1443.000000000,279.08
1444.000000000,0.0000
1445.000000000,0.0000
1446.000000000,52.603
1447.000000000,0.0000
1448.000000000,0.0000
1449.000000000,0.0000
1450.000000000,0.0000
1451.000000000,0.0000
1452.000000000,269.63
1453.000000000,0.0000
1454.000000000,479.50
1455.000000000,0.74474
1456.000000000,0.0000
1457.000000000,0.0000
1458.000000000,0.0000
1459.000000000,0.0000
1460.000000000,118.88
1461.000000000,18.880
1462.000000000,3.0021
1463.000000000,287.82
1464.000000000,0.0000
1465.000000000,0.0000
1466.000000000,0.0000
1467.000000000,0.0000
1468.000000000,0.0000
1469.000000000,0.0000
1470.000000000,0.0000
1471.000000000,0.0000
1472.000000000,0.0000
1473.000000000,0.0000
1474.000000000,0.0000
1475.000000000,442.96
1476.000000000,876.60
1477.000000000,1928.7
1478.000000000,0.0000
1479.000000000,2462.7
1480.000000000,0.0000
1481.000000000,0.0000
1482.000000000,0.0000
1483.000000000,0.10956E-01
1484.000000000,0.0000
1485.000000000,0.0000
1486.000000000,0.0000
1487.000000000,0.0000
1488.000000000,0.0000
1489.000000000,140.30
1490.000000000,0.0000
1491.000000000,0.0000
1492.000000000,0.0000
1493.000000000,0.0000
1494.000000000,0.0000
1495.000000000,0.0000
1496.000000000,1.1768
1497.000000000,77.480
1498.000000000,0.0000
1499.000000000,0.0000
1500.000000000,0.0000
1501.000000000,0.0000
1502.000000000,0.0000
1503.000000000,0.0000
1504.000000000,0.0000
1505.000000000,2.7095
1506.000000000,7950.9
1507.000000000,0.0000
1508.000000000,0.0000
1509.000000000,146.74
1510.000000000,0.0000
1511.000000000,0.0000
1512.000000000,1050.3
1513.000000000,0.0000
1514.000000000,0.0000
1515.000000000,0.0000
1516.000000000,0.0000
1517.000000000,0.0000
1518.000000000,0.0000
1519.000000000,0.0000
1520.000000000,0.0000
1521.000000000,0.0000
1522.000000000,0.0000
1523.000000000,0.0000
1524.000000000,0.0000
1525.000000000,540.12
1526.000000000,0.0000
1527.000000000,0.0000
1528.000000000,0.0000
1529.000000000,0.0000
1530.000000000,0.0000
1531.000000000,135.89
1532.000000000,5.3138
1533.000000000,0.0000
1534.000000000,9.3347
1535.000000000,0.0000
1536.000000000,0.0000
1537.000000000,0.0000
1538.000000000,0.0000
1539.000000000,0.0000
1540.000000000,0.0000
1541.000000000,0.0000
1542.000000000,0.0000
1543.000000000,0.0000
1544.000000000,94.761
1545.000000000,0.0000
1546.000000000,0.0000
1547.000000000,0.0000
1548.000000000,0.0000
1549.000000000,3518.1
1550.000000000,0.0000
1551.000000000,0.0000
1552.000000000,0.0000
1553.000000000,6708.8
1554.000000000,0.0000
1555.000000000,0.0000
1556.000000000,0.0000
1557.000000000,0.0000
1558.000000000,0.0000
1559.000000000,0.0000
1560.000000000,0.0000
1561.000000000,0.0000
1562.000000000,2177.6
1563.000000000,603.83
1564.000000000,705.68
1565.000000000,2995.6
1566.000000000,0.0000
1567.000000000,205.99
1568.000000000,1017.9
1569.000000000,0.0000
1570.000000000,0.0000
1571.000000000,0.0000
1572.000000000,0.0000
1573.000000000,0.0000
1574.000000000,0.0000
1575.000000000,0.0000
1576.000000000,0.0000
1577.000000000,0.0000
1578.000000000,0.0000
1579.000000000,0.0000
1580.000000000,0.0000
1581.000000000,0.0000
1582.000000000,0.0000
1583.000000000,0.0000
1584.000000000,0.0000
1585.000000000,0.0000
1586.000000000,0.0000
1587.000000000,0.0000
1588.000000000,0.0000
1589.000000000,0.0000
1590.000000000,2.7980
1591.000000000,0.0000
1592.000000000,2778.2
1593.000000000,0.0000
1594.000000000,0.0000
1595.000000000,0.0000
1596.000000000,0.0000
1597.000000000,0.0000
1598.000000000,68.404
1599.000000000,0.0000
1600.000000000,0.0000
1601.000000000,5443.4
1602.000000000,357.90
1603.000000000,4499.6
1604.000000000,52.226
1605.000000000,161.93
1606.000000000,0.0000
1607.000000000,0.0000
1608.000000000,0.0000
1609.000000000,0.0000
1610.000000000,5474.8
1611.000000000,97.526
1612.000000000,17869.
1613.000000000,2067.5
1614.000000000,433.01
1615.000000000,1230.8
1616.000000000,3087.6
1617.000000000,402.93
1618.000000000,0.0000
1619.000000000,0.0000
1620.000000000,0.0000
1621.000000000,0.0000
1622.000000000,0.0000
1623.000000000,0.0000
1624.000000000,0.0000
1625.000000000,0.0000
1626.000000000,0.0000
1627.000000000,0.0000
1628.000000000,27.984
1629.000000000,0.12529
1630.000000000,0.0000
1631.000000000,0.0000
1632.000000000,0.0000
1633.000000000,0.0000
1634.000000000,0.0000
1635.000000000,0.0000
1636.000000000,67.892
1637.000000000,0.0000
1638.000000000,41.818
1639.000000000,1498.2
1640.000000000,294.98
1641.000000000,0.0000
1642.000000000,0.0000
1643.000000000,0.0000
1644.000000000,11.281
1645.000000000,0.0000
1646.000000000,0.0000
1647.000000000,176.00
1648.000000000,228.21
1649.000000000,2091.0
1650.000000000,2618.2
1651.000000000,0.0000
1652.000000000,0.0000
1653.000000000,0.0000
1654.000000000,0.0000
1655.000000000,29.762
1656.000000000,439.50
1657.000000000,947.46
1658.000000000,1484.2
1659.000000000,698.90
1660.000000000,312.74
1661.000000000,256.58
1662.000000000,0.0000
1663.000000000,0.0000
1664.000000000,0.0000
1665.000000000,20.166
1666.000000000,5212.2
1667.000000000,40.973
1668.000000000,0.0000
1669.000000000,0.0000
1670.000000000,0.0000
1671.000000000,0.0000
1672.000000000,0.0000
1673.000000000,625.71
1674.000000000,300.34
1675.000000000,888.93
1676.000000000,1023.0
1677.000000000,0.0000
1678.000000000,82.814
1679.000000000,0.52773
1680.000000000,0.99109E-01
1681.000000000,321.69
1682.000000000,6721.5
1683.000000000,2.2540
1684.000000000,64.568
1685.000000000,0.0000
1686.000000000,0.0000
1687.000000000,1.0446
1688.000000000,0.65330E-01
1689.000000000,480.08
1690.000000000,229.62
1691.000000000,0.0000
1692.000000000,15.840
1693.000000000,0.0000
1694.000000000,0.0000
1695.000000000,0.0000
1696.000000000,4.7885
1697.000000000,1648.3
1698.000000000,2014.1
1699.000000000,247.99
1700.000000000,1262.8
1701.000000000,18.961
1702.000000000,0.0000
1703.000000000,0.0000
1704.000000000,0.0000
1705.000000000,0.0000
1706.000000000,0.0000
1707.000000000,0.0000
1708.000000000,78.583
1709.000000000,0.0000
1710.000000000,34.049
1711.000000000,0.0000
1712.000000000,0.0000
1713.000000000,0.0000
1714.000000000,0.0000
1715.000000000,0.0000
1716.000000000,0.0000
1717.000000000,0.0000
1718.000000000,0.0000
1719.000000000,0.0000
1720.000000000,0.0000
1721.000000000,0.0000
1722.000000000,0.0000
1723.000000000,0.0000
1724.000000000,124.38
1725.000000000,0.0000
1726.000000000,0.0000
1727.000000000,100.00
1728.000000000,0.0000
1729.000000000,5866.1
1730.000000000,3461.8
1731.000000000,11792.
1732.000000000,11616.
1733.000000000,5222.2
1734.000000000,1634.3
1735.000000000,567.76
1736.000000000,0.0000
1737.000000000,0.0000
1738.000000000,3422.1
1739.000000000,564.00
1740.000000000,0.0000
1741.000000000,0.0000
1742.000000000,0.0000
1743.000000000,0.0000
1744.000000000,1800.2
1745.000000000,101.10
1746.000000000,0.0000
1747.000000000,0.0000
1748.000000000,0.0000
1749.000000000,0.0000
1750.000000000,31.964
1751.000000000,0.0000
1752.000000000,0.0000
1753.000000000,0.0000
1754.000000000,0.0000
1755.000000000,0.0000
1756.000000000,0.0000
1757.000000000,0.0000
1758.000000000,0.0000
1759.000000000,0.0000
1760.000000000,0.0000
1761.000000000,0.0000
1762.000000000,0.0000
1763.000000000,0.0000
1764.000000000,0.0000
1765.000000000,0.0000
1766.000000000,30.707
1767.000000000,0.0000
1768.000000000,0.0000
1769.000000000,0.0000
1770.000000000,0.0000
1771.000000000,0.0000
1772.000000000,0.0000
1773.000000000,0.0000
1774.000000000,68.646
1775.000000000,0.0000
1776.000000000,0.0000
1777.000000000,537.74
1778.000000000,0.23949E-02
1779.000000000,151.06
1780.000000000,0.0000
1781.000000000,0.0000
1782.000000000,0.0000
1783.000000000,0.0000
1784.000000000,0.0000
1785.000000000,0.0000
1786.000000000,0.0000
1787.000000000,0.0000
1788.000000000,0.0000
1789.000000000,0.0000
1790.000000000,0.0000
1791.000000000,0.0000
1792.000000000,0.0000
1793.000000000,0.0000
1794.000000000,0.0000
1795.000000000,0.0000
1796.000000000,0.0000
1797.000000000,0.0000
1798.000000000,0.0000
1799.000000000,0.0000
1800.000000000,0.0000
1801.000000000,1571.9
1802.000000000,5761.5
1803.000000000,1595.0
1804.000000000,0.0000
1805.000000000,0.0000
1806.000000000,0.0000
1807.000000000,0.0000
1808.000000000,0.0000
1809.000000000,0.0000
1810.000000000,0.0000
1811.000000000,223.44
1812.000000000,2041.0
1813.000000000,0.66706E-02
1814.000000000,411.54
1815.000000000,16.976
1816.000000000,0.0000
1817.000000000,0.0000
1818.000000000,55.755
1819.000000000,0.0000
1820.000000000,0.0000
1821.000000000,0.0000
1822.000000000,224.29
1823.000000000,117.32
1824.000000000,0.60518
1825.000000000,30.617
1826.000000000,0.0000
1827.000000000,0.0000
1828.000000000,63.253
1829.000000000,0.0000
1830.000000000,0.0000
1831.000000000,0.13577
1832.000000000,0.0000
1833.000000000,0.0000
1834.000000000,0.0000
1835.000000000,0.0000
1836.000000000,0.0000
1837.000000000,0.0000
1838.000000000,0.0000
1839.000000000,0.0000
1840.000000000,0.0000
1841.000000000,0.0000
1842.000000000,109.10
1843.000000000,0.0000
1844.000000000,0.0000
1845.000000000,92.575
1846.000000000,59.459
1847.000000000,0.0000
1848.000000000,0.0000
1849.000000000,0.0000
1850.000000000,0.0000
1851.000000000,0.0000
1852.000000000,0.0000
1853.000000000,0.0000
1854.000000000,0.0000
1855.000000000,0.0000
1856.000000000,0.0000
1857.000000000,0.0000
1858.000000000,0.0000
1859.000000000,0.0000
1860.000000000,122.47
1861.000000000,0.0000
1862.000000000,0.0000
1863.000000000,0.0000
1864.000000000,55.095
1865.000000000,0.0000
1866.000000000,0.0000
1867.000000000,0.10519
1868.000000000,0.0000
1869.000000000,0.0000
1870.000000000,390.36
1871.000000000,133.64
1872.000000000,0.0000
1873.000000000,0.0000
1874.000000000,0.0000
1875.000000000,1.6487
1876.000000000,576.70
1877.000000000,1660.1
1878.000000000,6667.7
1879.000000000,484.91
1880.000000000,22.870
1881.000000000,143.90
1882.000000000,0.0000
1883.000000000,0.0000
1884.000000000,0.0000
1885.000000000,0.41617
1886.000000000,346.04
1887.000000000,0.0000
1888.000000000,0.0000
1889.000000000,0.0000
1890.000000000,0.0000
1891.000000000,0.0000
1892.000000000,0.0000
1893.000000000,0.0000
1894.000000000,0.0000
1895.000000000,0.0000
1896.000000000,0.0000
1897.000000000,0.0000
1898.000000000,0.0000
1899.000000000,0.0000
1900.000000000,0.0000
1901.000000000,0.0000
1902.000000000,0.0000
1903.000000000,0.0000
1904.000000000,0.0000
1905.000000000,0.0000
1906.000000000,0.0000
1907.000000000,0.0000
1908.000000000,0.0000
1909.000000000,0.0000
1910.000000000,0.0000
1911.000000000,0.0000
1912.000000000,0.0000
1913.000000000,327.86
1914.000000000,0.0000
1915.000000000,0.0000
1916.000000000,0.0000
1917.000000000,0.0000
1918.000000000,0.0000
1919.000000000,0.0000
1920.000000000,0.0000
1921.000000000,0.0000
1922.000000000,0.0000
1923.000000000,0.0000
1924.000000000,0.0000
1925.000000000,0.0000
1926.000000000,0.0000
1927.000000000,0.0000
1928.000000000,0.0000
1929.000000000,0.0000
1930.000000000,177.20
1931.000000000,0.0000
1932.000000000,0.0000
1933.000000000,0.0000
1934.000000000,0.0000
1935.000000000,0.0000
1936.000000000,0.0000
1937.000000000,27.029
1938.000000000,106.99
1939.000000000,0.0000
1940.000000000,0.0000
1941.000000000,0.0000
1942.000000000,1095.9
1943.000000000,0.0000
1944.000000000,0.0000
1945.000000000,0.0000
1946.000000000,0.0000
1947.000000000,0.0000
1948.000000000,0.0000
1949.000000000,337.13
1950.000000000,7647.3
1951.000000000,1202.9
1952.000000000,0.0000
1953.000000000,0.0000
1954.000000000,0.0000
1955.000000000,0.0000
1956.000000000,0.0000
1957.000000000,0.0000
1958.000000000,0.0000
1959.000000000,0.0000
1960.000000000,0.0000
1961.000000000,0.0000
1962.000000000,0.0000
1963.000000000,0.0000
1964.000000000,56.812
1965.000000000,3.1257
1966.000000000,705.69
1967.000000000,7333.7
1968.000000000,168.34
1969.000000000,0.0000
1970.000000000,0.0000
1971.000000000,0.0000
1972.000000000,0.0000
1973.000000000,0.0000
1974.000000000,0.0000
1975.000000000,0.0000
1976.000000000,0.0000
1977.000000000,0.0000
1978.000000000,0.0000
1979.000000000,0.0000
1980.000000000,0.0000
1981.000000000,385.20
1982.000000000,0.0000
1983.000000000,0.0000
1984.000000000,0.0000
1985.000000000,0.0000
1986.000000000,0.0000
1987.000000000,0.0000
1988.000000000,16.108
1989.000000000,0.0000
1990.000000000,0.0000
1991.000000000,1.9794
1992.000000000,0.0000
1993.000000000,0.0000
1994.000000000,0.0000
1995.000000000,29.415
1996.000000000,505.58
1997.000000000,0.39436
1998.000000000,0.0000
1999.000000000,101.15
2000.000000000,0.0000
2001.000000000,0.0000
2002.000000000,0.0000
2003.000000000,0.0000
2004.000000000,7.6978
2005.000000000,0.0000
2006.000000000,0.0000
2007.000000000,425.54
2008.000000000,0.0000
2009.000000000,0.0000
2010.000000000,0.0000
2011.000000000,0.0000
2012.000000000,771.11
2013.000000000,1340.1
2014.000000000,3129.3
2015.000000000,3304.6
2016.000000000,1401.6
2017.000000000,2320.1
2018.000000000,0.0000
2019.000000000,0.0000
2020.000000000,0.0000
2021.000000000,0.0000
2022.000000000,0.0000
2023.000000000,0.0000
2024.000000000,0.0000
2025.000000000,0.0000
2026.000000000,0.0000
2027.000000000,0.0000
2028.000000000,0.0000
2029.000000000,0.0000
2030.000000000,0.0000
2031.000000000,0.0000
2032.000000000,0.0000
2033.000000000,0.18818E-01
2034.000000000,0.0000
2035.000000000,0.0000
2036.000000000,0.0000
2037.000000000,0.0000
2038.000000000,7534.3
2039.000000000,214.46
2040.000000000,0.0000
2041.000000000,0.0000
2042.000000000,0.0000
2043.000000000,0.0000
2044.000000000,0.0000
2045.000000000,0.0000
2046.000000000,0.0000
2047.000000000,0.0000
2048.000000000,33.800
2049.000000000,2860.4
2050.000000000,1990.1
2051.000000000,2634.4
2052.000000000,635.19
2053.000000000,0.0000
2054.000000000,0.0000
2055.000000000,0.0000
2056.000000000,0.0000
2057.000000000,0.0000
2058.000000000,625.47
2059.000000000,1201.7
2060.000000000,0.0000
2061.000000000,0.0000
2062.000000000,0.0000
2063.000000000,0.0000
2064.000000000,0.0000
2065.000000000,0.0000
2066.000000000,0.0000
2067.000000000,0.0000
2068.000000000,0.0000
2069.000000000,0.0000
