time,SOUTHOUT
1.000000000000,-183.18
2.000000000000,-183.19
3.000000000000,-183.28
4.000000000000,-183.98
5.000000000000,-184.09
6.000000000000,-183.97
7.000000000000,-184.04
8.000000000000,-184.17
9.000000000000,-187.67
10.00000000000,-189.68
11.00000000000,-186.87
12.00000000000,-186.09
13.00000000000,-185.71
14.00000000000,-185.54
15.00000000000,-185.49
16.00000000000,-185.47
17.00000000000,-185.49
18.00000000000,-185.52
19.00000000000,-185.58
20.00000000000,-185.63
21.00000000000,-185.70
22.00000000000,-185.76
23.00000000000,-185.81
24.00000000000,-185.85
25.00000000000,-185.88
26.00000000000,-185.92
27.00000000000,-185.95
28.00000000000,-185.99
29.00000000000,-186.02
30.00000000000,-186.05
31.00000000000,-186.09
32.00000000000,-186.12
33.00000000000,-186.14
34.00000000000,-186.17
35.00000000000,-186.20
36.00000000000,-186.22
37.00000000000,-186.25
38.00000000000,-186.27
39.00000000000,-186.29
40.00000000000,-186.32
41.00000000000,-186.36
42.00000000000,-186.36
43.00000000000,-186.36
44.00000000000,-186.36
45.00000000000,-186.36
46.00000000000,-186.36
47.00000000000,-186.36
48.00000000000,-186.36
49.00000000000,-186.36
50.00000000000,-186.36
51.00000000000,-186.36
52.00000000000,-186.55
53.00000000000,-186.43
54.00000000000,-186.40
55.00000000000,-186.38
56.00000000000,-186.55
57.00000000000,-186.43
58.00000000000,-186.40
59.00000000000,-186.37
60.00000000000,-186.36
61.00000000000,-186.35
62.00000000000,-186.34
63.00000000000,-186.34
64.00000000000,-186.33
65.00000000000,-186.33
66.00000000000,-186.33
67.00000000000,-186.32
68.00000000000,-186.32
69.00000000000,-186.90
70.00000000000,-186.54
71.00000000000,-186.45
72.00000000000,-186.40
73.00000000000,-186.37
74.00000000000,-186.36
75.00000000000,-186.34
76.00000000000,-186.34
77.00000000000,-186.33
78.00000000000,-186.32
79.00000000000,-186.32
80.00000000000,-186.32
81.00000000000,-186.31
82.00000000000,-186.64
83.00000000000,-186.44
84.00000000000,-186.38
85.00000000000,-186.35
86.00000000000,-186.33
87.00000000000,-186.32
88.00000000000,-186.31
89.00000000000,-186.31
90.00000000000,-186.31
91.00000000000,-186.30
92.00000000000,-186.30
93.00000000000,-187.75
94.00000000000,-186.88
95.00000000000,-186.62
96.00000000000,-186.49
97.00000000000,-186.41
98.00000000000,-186.36
99.00000000000,-186.33
100.0000000000,-186.31
101.0000000000,-186.29
102.0000000000,-186.28
103.0000000000,-186.27
104.0000000000,-186.26
105.0000000000,-186.26
106.0000000000,-186.25
107.0000000000,-186.25
108.0000000000,-187.08
109.0000000000,-186.56
110.0000000000,-186.42
111.0000000000,-186.34
112.0000000000,-186.30
113.0000000000,-186.27
114.0000000000,-186.25
115.0000000000,-186.23
116.0000000000,-186.22
117.0000000000,-186.21
118.0000000000,-188.95
119.0000000000,-191.94
120.0000000000,-188.62
121.0000000000,-187.62
122.0000000000,-188.83
123.0000000000,-187.43
124.0000000000,-186.94
125.0000000000,-186.66
126.0000000000,-186.49
127.0000000000,-186.38
128.0000000000,-186.31
129.0000000000,-186.25
130.0000000000,-187.11
131.0000000000,-187.64
132.0000000000,-186.79
133.0000000000,-186.52
134.0000000000,-186.36
135.0000000000,-187.72
136.0000000000,-186.76
137.0000000000,-186.48
138.0000000000,-186.33
139.0000000000,-186.23
140.0000000000,-186.17
141.0000000000,-186.13
142.0000000000,-186.09
143.0000000000,-186.07
144.0000000000,-189.33
145.0000000000,-187.57
146.0000000000,-191.97
147.0000000000,-188.50
148.0000000000,-187.47
149.0000000000,-187.62
150.0000000000,-186.86
151.0000000000,-186.54
152.0000000000,-186.34
153.0000000000,-186.22
154.0000000000,-186.25
155.0000000000,-186.13
156.0000000000,-186.07
157.0000000000,-186.03
158.0000000000,-186.03
159.0000000000,-187.15
160.0000000000,-186.42
161.0000000000,-186.22
162.0000000000,-186.10
163.0000000000,-186.03
164.0000000000,-185.98
165.0000000000,-186.68
166.0000000000,-192.77
167.0000000000,-189.10
168.0000000000,-187.66
169.0000000000,-187.45
170.0000000000,-186.90
171.0000000000,-186.49
172.0000000000,-186.27
173.0000000000,-186.13
174.0000000000,-186.04
175.0000000000,-185.98
176.0000000000,-185.94
177.0000000000,-185.91
178.0000000000,-185.89
179.0000000000,-185.87
180.0000000000,-185.85
181.0000000000,-187.47
182.0000000000,-186.47
183.0000000000,-186.55
184.0000000000,-186.18
185.0000000000,-186.03
186.0000000000,-185.94
187.0000000000,-185.88
188.0000000000,-185.84
189.0000000000,-185.81
190.0000000000,-185.79
191.0000000000,-185.77
192.0000000000,-185.76
193.0000000000,-185.75
194.0000000000,-185.74
195.0000000000,-185.73
196.0000000000,-186.13
197.0000000000,-190.15
198.0000000000,-189.71
199.0000000000,-188.01
200.0000000000,-187.67
201.0000000000,-186.77
202.0000000000,-186.48
203.0000000000,-186.35
204.0000000000,-186.07
205.0000000000,-185.94
206.0000000000,-185.85
207.0000000000,-185.80
208.0000000000,-185.95
209.0000000000,-185.80
210.0000000000,-186.38
211.0000000000,-185.96
212.0000000000,-185.84
213.0000000000,-185.76
214.0000000000,-185.72
215.0000000000,-185.69
216.0000000000,-185.66
217.0000000000,-185.65
218.0000000000,-185.63
219.0000000000,-185.62
220.0000000000,-185.61
221.0000000000,-185.60
222.0000000000,-185.59
223.0000000000,-185.62
224.0000000000,-185.80
225.0000000000,-185.66
226.0000000000,-185.62
227.0000000000,-185.59
228.0000000000,-185.57
229.0000000000,-185.56
230.0000000000,-185.55
231.0000000000,-185.54
232.0000000000,-185.53
233.0000000000,-185.52
234.0000000000,-185.64
235.0000000000,-185.56
236.0000000000,-188.96
237.0000000000,-186.92
238.0000000000,-186.80
239.0000000000,-190.60
240.0000000000,-191.21
241.0000000000,-188.13
242.0000000000,-187.07
243.0000000000,-186.48
244.0000000000,-186.13
245.0000000000,-185.92
246.0000000000,-187.33
247.0000000000,-186.29
248.0000000000,-187.19
249.0000000000,-187.01
250.0000000000,-186.25
251.0000000000,-185.96
252.0000000000,-186.77
253.0000000000,-186.23
254.0000000000,-186.40
255.0000000000,-185.94
256.0000000000,-185.77
257.0000000000,-185.66
258.0000000000,-185.60
259.0000000000,-185.55
260.0000000000,-186.36
261.0000000000,-187.46
262.0000000000,-186.69
263.0000000000,-195.87
264.0000000000,-197.57
265.0000000000,-190.96
266.0000000000,-188.73
267.0000000000,-187.50
268.0000000000,-186.78
269.0000000000,-186.35
270.0000000000,-186.08
271.0000000000,-185.90
272.0000000000,-187.11
273.0000000000,-186.22
274.0000000000,-185.95
275.0000000000,-185.80
276.0000000000,-185.71
277.0000000000,-185.64
278.0000000000,-185.60
279.0000000000,-185.58
280.0000000000,-185.55
281.0000000000,-185.54
282.0000000000,-185.52
283.0000000000,-185.51
284.0000000000,-185.50
285.0000000000,-185.49
286.0000000000,-185.52
287.0000000000,-186.68
288.0000000000,-188.10
289.0000000000,-193.16
290.0000000000,-188.82
291.0000000000,-187.40
292.0000000000,-186.69
293.0000000000,-186.24
294.0000000000,-185.97
295.0000000000,-185.80
296.0000000000,-185.70
297.0000000000,-185.63
298.0000000000,-185.58
299.0000000000,-185.54
300.0000000000,-185.52
301.0000000000,-185.50
302.0000000000,-185.48
303.0000000000,-185.47
304.0000000000,-185.51
305.0000000000,-185.47
306.0000000000,-185.45
307.0000000000,-185.44
308.0000000000,-186.28
309.0000000000,-185.99
310.0000000000,-186.42
311.0000000000,-186.45
312.0000000000,-185.91
313.0000000000,-186.39
314.0000000000,-185.85
315.0000000000,-185.67
316.0000000000,-185.71
317.0000000000,-185.59
318.0000000000,-185.50
319.0000000000,-185.46
320.0000000000,-185.42
321.0000000000,-185.40
322.0000000000,-185.38
323.0000000000,-185.37
324.0000000000,-185.36
325.0000000000,-185.35
326.0000000000,-185.61
327.0000000000,-185.70
328.0000000000,-187.25
329.0000000000,-187.51
330.0000000000,-186.35
331.0000000000,-185.92
332.0000000000,-185.69
333.0000000000,-185.55
334.0000000000,-185.47
335.0000000000,-185.41
336.0000000000,-185.37
337.0000000000,-185.35
338.0000000000,-185.33
339.0000000000,-185.31
340.0000000000,-185.63
341.0000000000,-185.42
342.0000000000,-185.36
343.0000000000,-185.32
344.0000000000,-185.30
345.0000000000,-185.28
346.0000000000,-185.26
347.0000000000,-185.25
348.0000000000,-185.25
349.0000000000,-185.24
350.0000000000,-185.23
351.0000000000,-185.22
352.0000000000,-185.22
353.0000000000,-185.21
354.0000000000,-185.20
355.0000000000,-186.50
356.0000000000,-186.18
357.0000000000,-185.67
358.0000000000,-185.48
359.0000000000,-185.36
360.0000000000,-185.72
361.0000000000,-186.29
362.0000000000,-186.41
363.0000000000,-185.75
364.0000000000,-185.51
365.0000000000,-185.38
366.0000000000,-185.30
367.0000000000,-185.25
368.0000000000,-185.21
369.0000000000,-185.19
370.0000000000,-185.17
371.0000000000,-185.15
372.0000000000,-185.14
373.0000000000,-185.13
374.0000000000,-185.13
375.0000000000,-185.12
376.0000000000,-185.11
377.0000000000,-185.10
378.0000000000,-185.10
379.0000000000,-185.09
380.0000000000,-185.09
381.0000000000,-185.08
382.0000000000,-185.07
383.0000000000,-185.07
384.0000000000,-185.06
385.0000000000,-185.06
386.0000000000,-185.05
387.0000000000,-185.05
388.0000000000,-185.04
389.0000000000,-185.15
390.0000000000,-185.08
391.0000000000,-185.06
392.0000000000,-185.04
393.0000000000,-185.03
394.0000000000,-185.02
395.0000000000,-185.01
396.0000000000,-185.01
397.0000000000,-185.00
398.0000000000,-184.99
399.0000000000,-184.99
400.0000000000,-184.98
401.0000000000,-184.98
402.0000000000,-184.97
403.0000000000,-184.97
404.0000000000,-184.96
405.0000000000,-184.96
406.0000000000,-184.95
407.0000000000,-184.95
408.0000000000,-184.94
409.0000000000,-184.94
410.0000000000,-184.93
411.0000000000,-184.93
412.0000000000,-184.92
413.0000000000,-184.92
414.0000000000,-184.91
415.0000000000,-184.91
416.0000000000,-184.90
417.0000000000,-184.90
418.0000000000,-184.89
419.0000000000,-184.89
420.0000000000,-184.88
421.0000000000,-184.96
422.0000000000,-186.03
423.0000000000,-185.67
424.0000000000,-185.27
425.0000000000,-185.11
426.0000000000,-185.05
427.0000000000,-184.97
428.0000000000,-184.93
429.0000000000,-184.90
430.0000000000,-184.88
431.0000000000,-184.87
432.0000000000,-184.85
433.0000000000,-184.85
434.0000000000,-184.89
435.0000000000,-184.85
436.0000000000,-184.84
437.0000000000,-184.83
438.0000000000,-184.82
439.0000000000,-184.81
440.0000000000,-184.81
441.0000000000,-184.80
442.0000000000,-184.80
443.0000000000,-184.79
444.0000000000,-184.79
445.0000000000,-184.79
446.0000000000,-184.78
447.0000000000,-184.78
448.0000000000,-185.03
449.0000000000,-184.87
450.0000000000,-184.83
451.0000000000,-184.85
452.0000000000,-184.81
453.0000000000,-184.79
454.0000000000,-184.78
455.0000000000,-184.77
456.0000000000,-184.76
457.0000000000,-184.76
458.0000000000,-184.75
459.0000000000,-185.70
460.0000000000,-185.11
461.0000000000,-185.00
462.0000000000,-184.90
463.0000000000,-184.94
464.0000000000,-184.84
465.0000000000,-184.80
466.0000000000,-184.77
467.0000000000,-184.76
468.0000000000,-184.74
469.0000000000,-184.75
470.0000000000,-184.73
471.0000000000,-184.72
472.0000000000,-184.72
473.0000000000,-184.71
474.0000000000,-184.70
475.0000000000,-184.82
476.0000000000,-184.75
477.0000000000,-184.72
478.0000000000,-184.71
479.0000000000,-184.70
480.0000000000,-184.69
481.0000000000,-184.69
482.0000000000,-184.68
483.0000000000,-184.68
484.0000000000,-184.67
485.0000000000,-184.67
486.0000000000,-184.66
487.0000000000,-184.66
488.0000000000,-184.66
489.0000000000,-184.65
490.0000000000,-184.65
491.0000000000,-184.65
492.0000000000,-185.37
493.0000000000,-184.92
494.0000000000,-185.13
495.0000000000,-185.50
496.0000000000,-185.02
497.0000000000,-184.89
498.0000000000,-185.49
499.0000000000,-185.16
500.0000000000,-184.91
501.0000000000,-184.80
502.0000000000,-184.74
503.0000000000,-184.70
504.0000000000,-184.67
505.0000000000,-184.65
506.0000000000,-184.63
507.0000000000,-184.62
508.0000000000,-184.89
509.0000000000,-184.73
510.0000000000,-185.36
511.0000000000,-189.49
512.0000000000,-186.84
513.0000000000,-185.85
514.0000000000,-185.36
515.0000000000,-185.08
516.0000000000,-184.91
517.0000000000,-184.81
518.0000000000,-184.74
519.0000000000,-184.70
520.0000000000,-184.67
521.0000000000,-184.65
522.0000000000,-184.63
523.0000000000,-184.62
524.0000000000,-184.61
525.0000000000,-184.67
526.0000000000,-184.67
527.0000000000,-184.63
528.0000000000,-184.75
529.0000000000,-185.59
530.0000000000,-186.71
531.0000000000,-185.50
532.0000000000,-185.11
533.0000000000,-184.90
534.0000000000,-184.78
535.0000000000,-184.70
536.0000000000,-194.72
537.0000000000,-192.76
538.0000000000,-189.91
539.0000000000,-187.47
540.0000000000,-186.45
541.0000000000,-189.43
542.0000000000,-186.78
543.0000000000,-185.94
544.0000000000,-185.52
545.0000000000,-185.21
546.0000000000,-185.03
547.0000000000,-184.91
548.0000000000,-184.83
549.0000000000,-184.79
550.0000000000,-184.75
551.0000000000,-184.72
552.0000000000,-184.70
553.0000000000,-184.68
554.0000000000,-184.67
555.0000000000,-184.66
556.0000000000,-184.69
557.0000000000,-184.71
558.0000000000,-185.43
559.0000000000,-184.94
560.0000000000,-184.80
561.0000000000,-184.73
562.0000000000,-185.68
563.0000000000,-186.24
564.0000000000,-186.21
565.0000000000,-185.36
566.0000000000,-185.05
567.0000000000,-184.87
568.0000000000,-184.77
569.0000000000,-184.70
570.0000000000,-184.66
571.0000000000,-185.05
572.0000000000,-184.77
573.0000000000,-184.68
574.0000000000,-184.63
575.0000000000,-184.60
576.0000000000,-184.58
577.0000000000,-184.56
578.0000000000,-184.55
579.0000000000,-186.32
580.0000000000,-189.89
581.0000000000,-186.72
582.0000000000,-185.81
583.0000000000,-185.31
584.0000000000,-185.02
585.0000000000,-184.84
586.0000000000,-184.73
587.0000000000,-184.66
588.0000000000,-184.61
589.0000000000,-185.06
590.0000000000,-185.87
591.0000000000,-185.09
592.0000000000,-184.85
593.0000000000,-184.71
594.0000000000,-184.92
595.0000000000,-186.12
596.0000000000,-186.93
597.0000000000,-185.57
598.0000000000,-185.13
599.0000000000,-184.88
600.0000000000,-184.74
601.0000000000,-184.65
602.0000000000,-184.59
603.0000000000,-184.55
604.0000000000,-184.52
605.0000000000,-184.54
606.0000000000,-184.50
607.0000000000,-184.70
608.0000000000,-184.61
609.0000000000,-184.53
610.0000000000,-184.49
611.0000000000,-184.47
612.0000000000,-184.48
613.0000000000,-185.87
614.0000000000,-185.39
615.0000000000,-184.91
616.0000000000,-185.76
617.0000000000,-185.01
618.0000000000,-184.76
619.0000000000,-184.63
620.0000000000,-184.58
621.0000000000,-184.92
622.0000000000,-184.95
623.0000000000,-184.69
624.0000000000,-184.56
625.0000000000,-184.74
626.0000000000,-184.55
627.0000000000,-186.96
628.0000000000,-185.62
629.0000000000,-186.27
630.0000000000,-185.98
631.0000000000,-185.18
632.0000000000,-184.87
633.0000000000,-184.71
634.0000000000,-184.65
635.0000000000,-189.95
636.0000000000,-187.52
637.0000000000,-186.02
638.0000000000,-185.37
639.0000000000,-185.00
640.0000000000,-184.78
641.0000000000,-184.64
642.0000000000,-184.55
643.0000000000,-184.49
644.0000000000,-184.45
645.0000000000,-184.42
646.0000000000,-184.40
647.0000000000,-184.38
648.0000000000,-184.37
649.0000000000,-186.61
650.0000000000,-185.22
651.0000000000,-184.85
652.0000000000,-184.65
653.0000000000,-184.53
654.0000000000,-184.46
655.0000000000,-184.41
656.0000000000,-184.38
657.0000000000,-184.36
658.0000000000,-184.34
659.0000000000,-184.42
660.0000000000,-184.78
661.0000000000,-185.78
662.0000000000,-184.91
663.0000000000,-184.66
664.0000000000,-184.51
665.0000000000,-184.43
666.0000000000,-184.38
667.0000000000,-184.34
668.0000000000,-184.32
669.0000000000,-184.30
670.0000000000,-184.29
671.0000000000,-184.28
672.0000000000,-184.27
673.0000000000,-184.26
674.0000000000,-191.80
675.0000000000,-191.34
676.0000000000,-187.69
677.0000000000,-186.37
678.0000000000,-185.55
679.0000000000,-185.09
680.0000000000,-184.81
681.0000000000,-184.64
682.0000000000,-184.52
683.0000000000,-184.45
684.0000000000,-184.40
685.0000000000,-184.36
686.0000000000,-184.33
687.0000000000,-184.31
688.0000000000,-184.30
689.0000000000,-184.29
690.0000000000,-184.28
691.0000000000,-184.27
692.0000000000,-184.94
693.0000000000,-184.52
694.0000000000,-184.40
695.0000000000,-184.34
696.0000000000,-184.30
697.0000000000,-184.28
698.0000000000,-184.26
699.0000000000,-184.24
700.0000000000,-184.23
701.0000000000,-184.23
702.0000000000,-184.22
703.0000000000,-184.21
704.0000000000,-184.21
705.0000000000,-184.20
706.0000000000,-184.20
707.0000000000,-184.19
708.0000000000,-184.19
709.0000000000,-184.19
710.0000000000,-184.22
711.0000000000,-184.19
712.0000000000,-184.18
713.0000000000,-184.17
714.0000000000,-184.16
715.0000000000,-184.16
716.0000000000,-184.15
717.0000000000,-184.15
718.0000000000,-184.22
719.0000000000,-184.17
720.0000000000,-184.15
721.0000000000,-184.14
722.0000000000,-184.21
723.0000000000,-184.25
724.0000000000,-184.18
725.0000000000,-184.15
726.0000000000,-184.13
727.0000000000,-187.04
728.0000000000,-185.37
729.0000000000,-184.81
730.0000000000,-184.70
731.0000000000,-184.99
732.0000000000,-185.41
733.0000000000,-185.70
734.0000000000,-184.85
735.0000000000,-184.55
736.0000000000,-184.38
737.0000000000,-184.28
738.0000000000,-184.21
739.0000000000,-184.24
740.0000000000,-185.57
741.0000000000,-184.83
742.0000000000,-184.50
743.0000000000,-184.33
744.0000000000,-184.24
745.0000000000,-184.18
746.0000000000,-184.14
747.0000000000,-184.11
748.0000000000,-184.09
749.0000000000,-184.08
750.0000000000,-184.07
751.0000000000,-184.06
752.0000000000,-184.99
753.0000000000,-185.49
754.0000000000,-184.74
755.0000000000,-184.44
756.0000000000,-184.28
757.0000000000,-184.19
758.0000000000,-184.13
759.0000000000,-184.09
760.0000000000,-184.07
761.0000000000,-184.90
762.0000000000,-185.54
763.0000000000,-184.67
764.0000000000,-184.40
765.0000000000,-184.31
766.0000000000,-184.18
767.0000000000,-184.12
768.0000000000,-184.08
769.0000000000,-184.05
770.0000000000,-184.03
771.0000000000,-184.01
772.0000000000,-184.00
773.0000000000,-183.99
774.0000000000,-183.99
775.0000000000,-183.98
776.0000000000,-183.97
777.0000000000,-183.99
778.0000000000,-184.07
779.0000000000,-184.00
780.0000000000,-183.98
781.0000000000,-183.97
782.0000000000,-183.96
783.0000000000,-183.95
784.0000000000,-183.94
785.0000000000,-183.94
786.0000000000,-183.93
787.0000000000,-183.93
788.0000000000,-183.92
789.0000000000,-184.27
790.0000000000,-184.15
791.0000000000,-184.08
792.0000000000,-184.00
793.0000000000,-183.96
794.0000000000,-185.23
795.0000000000,-184.42
796.0000000000,-184.20
797.0000000000,-184.50
798.0000000000,-184.27
799.0000000000,-184.27
800.0000000000,-184.09
801.0000000000,-184.01
802.0000000000,-183.96
803.0000000000,-183.93
804.0000000000,-183.91
805.0000000000,-183.89
806.0000000000,-183.88
807.0000000000,-184.15
808.0000000000,-184.00
809.0000000000,-185.38
810.0000000000,-189.70
811.0000000000,-189.23
812.0000000000,-186.40
813.0000000000,-185.38
814.0000000000,-184.81
815.0000000000,-184.66
816.0000000000,-184.34
817.0000000000,-184.19
818.0000000000,-184.09
819.0000000000,-184.02
820.0000000000,-183.98
821.0000000000,-183.95
822.0000000000,-183.92
823.0000000000,-183.91
824.0000000000,-183.90
825.0000000000,-183.89
826.0000000000,-184.14
827.0000000000,-183.97
828.0000000000,-184.00
829.0000000000,-184.54
830.0000000000,-184.14
831.0000000000,-184.02
832.0000000000,-184.37
833.0000000000,-186.38
834.0000000000,-184.87
835.0000000000,-184.44
836.0000000000,-185.40
837.0000000000,-184.82
838.0000000000,-186.16
839.0000000000,-184.91
840.0000000000,-184.47
841.0000000000,-184.23
842.0000000000,-184.10
843.0000000000,-184.01
844.0000000000,-185.26
845.0000000000,-184.42
846.0000000000,-184.18
847.0000000000,-186.24
848.0000000000,-184.82
849.0000000000,-184.42
850.0000000000,-184.20
851.0000000000,-184.07
852.0000000000,-183.99
853.0000000000,-183.94
854.0000000000,-183.90
855.0000000000,-183.90
856.0000000000,-183.87
857.0000000000,-183.91
858.0000000000,-183.87
859.0000000000,-183.85
860.0000000000,-183.84
861.0000000000,-190.62
862.0000000000,-191.45
863.0000000000,-190.95
864.0000000000,-188.70
865.0000000000,-187.22
866.0000000000,-188.59
867.0000000000,-191.20
868.0000000000,-187.24
869.0000000000,-185.95
870.0000000000,-185.20
871.0000000000,-186.97
872.0000000000,-185.80
873.0000000000,-185.11
874.0000000000,-185.97
875.0000000000,-185.05
876.0000000000,-185.17
877.0000000000,-184.60
878.0000000000,-184.38
879.0000000000,-189.93
880.0000000000,-186.46
881.0000000000,-189.84
882.0000000000,-186.59
883.0000000000,-185.55
884.0000000000,-184.98
885.0000000000,-184.64
886.0000000000,-184.43
887.0000000000,-184.30
888.0000000000,-184.21
889.0000000000,-184.15
890.0000000000,-184.11
891.0000000000,-184.09
892.0000000000,-184.07
893.0000000000,-184.05
894.0000000000,-184.50
895.0000000000,-187.96
896.0000000000,-186.00
897.0000000000,-186.87
898.0000000000,-186.11
899.0000000000,-185.23
900.0000000000,-184.79
901.0000000000,-186.24
902.0000000000,-185.20
903.0000000000,-184.70
904.0000000000,-184.89
905.0000000000,-184.50
906.0000000000,-184.32
907.0000000000,-184.22
908.0000000000,-186.40
909.0000000000,-187.01
910.0000000000,-185.49
911.0000000000,-184.89
912.0000000000,-185.09
913.0000000000,-184.58
914.0000000000,-184.38
915.0000000000,-184.26
916.0000000000,-184.19
917.0000000000,-184.14
918.0000000000,-184.12
919.0000000000,-186.37
920.0000000000,-184.95
921.0000000000,-184.57
922.0000000000,-184.36
923.0000000000,-184.24
924.0000000000,-184.16
925.0000000000,-184.12
926.0000000000,-184.09
927.0000000000,-184.06
928.0000000000,-184.05
929.0000000000,-184.04
930.0000000000,-184.03
931.0000000000,-184.02
932.0000000000,-184.01
933.0000000000,-184.01
934.0000000000,-184.00
935.0000000000,-184.00
936.0000000000,-184.00
937.0000000000,-183.99
938.0000000000,-183.99
939.0000000000,-183.98
940.0000000000,-183.98
941.0000000000,-183.97
942.0000000000,-183.97
943.0000000000,-184.60
944.0000000000,-184.85
945.0000000000,-184.35
946.0000000000,-184.19
947.0000000000,-184.10
948.0000000000,-184.04
949.0000000000,-184.00
950.0000000000,-183.98
951.0000000000,-183.96
952.0000000000,-183.95
953.0000000000,-183.94
954.0000000000,-183.93
955.0000000000,-184.56
956.0000000000,-184.65
957.0000000000,-185.21
958.0000000000,-185.88
959.0000000000,-184.78
960.0000000000,-184.42
961.0000000000,-184.22
962.0000000000,-186.03
963.0000000000,-185.62
964.0000000000,-184.74
965.0000000000,-184.41
966.0000000000,-184.22
967.0000000000,-184.10
968.0000000000,-184.39
969.0000000000,-184.59
970.0000000000,-184.21
971.0000000000,-184.08
972.0000000000,-184.00
973.0000000000,-184.21
974.0000000000,-184.02
975.0000000000,-183.96
976.0000000000,-183.92
977.0000000000,-183.90
978.0000000000,-183.88
979.0000000000,-183.87
980.0000000000,-183.86
981.0000000000,-183.85
982.0000000000,-183.84
983.0000000000,-184.95
984.0000000000,-184.27
985.0000000000,-184.73
986.0000000000,-184.23
987.0000000000,-184.06
988.0000000000,-183.97
989.0000000000,-183.91
990.0000000000,-183.87
991.0000000000,-183.84
992.0000000000,-183.83
993.0000000000,-183.81
994.0000000000,-183.80
995.0000000000,-183.79
996.0000000000,-183.79
997.0000000000,-183.78
998.0000000000,-183.77
999.0000000000,-183.77
1000.000000000,-184.22
1001.000000000,-183.94
1002.000000000,-183.86
1003.000000000,-183.81
1004.000000000,-183.79
1005.000000000,-183.77
1006.000000000,-183.75
1007.000000000,-183.74
1008.000000000,-183.74
1009.000000000,-183.74
1010.000000000,-183.73
1011.000000000,-183.72
1012.000000000,-188.96
1013.000000000,-186.55
1014.000000000,-185.19
1015.000000000,-184.60
1016.000000000,-184.27
1017.000000000,-184.07
1018.000000000,-183.94
1019.000000000,-183.87
1020.000000000,-183.81
1021.000000000,-183.78
1022.000000000,-183.76
1023.000000000,-183.74
1024.000000000,-183.73
1025.000000000,-184.05
1026.000000000,-184.43
1027.000000000,-194.89
1028.000000000,-192.86
1029.000000000,-188.10
1030.000000000,-186.35
1031.000000000,-185.37
1032.000000000,-184.80
1033.000000000,-184.88
1034.000000000,-190.76
1035.000000000,-186.65
1036.000000000,-185.49
1037.000000000,-184.86
1038.000000000,-184.49
1039.000000000,-184.26
1040.000000000,-184.12
1041.000000000,-184.30
1042.000000000,-184.32
1043.000000000,-184.09
1044.000000000,-183.99
1045.000000000,-183.94
1046.000000000,-183.90
1047.000000000,-183.87
1048.000000000,-183.99
1049.000000000,-184.36
1050.000000000,-184.13
1051.000000000,-184.14
1052.000000000,-183.98
1053.000000000,-183.91
1054.000000000,-183.87
1055.000000000,-183.84
1056.000000000,-183.82
1057.000000000,-183.81
1058.000000000,-183.80
1059.000000000,-183.79
1060.000000000,-183.98
1061.000000000,-184.80
1062.000000000,-188.13
1063.000000000,-185.70
1064.000000000,-184.86
1065.000000000,-184.44
1066.000000000,-184.19
1067.000000000,-184.04
1068.000000000,-183.95
1069.000000000,-183.89
1070.000000000,-183.85
1071.000000000,-183.82
1072.000000000,-183.80
1073.000000000,-183.79
1074.000000000,-183.78
1075.000000000,-183.77
1076.000000000,-183.76
1077.000000000,-188.38
1078.000000000,-185.53
1079.000000000,-184.77
1080.000000000,-184.37
1081.000000000,-184.14
1082.000000000,-184.00
1083.000000000,-183.91
1084.000000000,-183.85
1085.000000000,-183.82
1086.000000000,-183.79
1087.000000000,-183.77
1088.000000000,-183.76
1089.000000000,-183.75
1090.000000000,-183.74
1091.000000000,-187.66
1092.000000000,-186.05
1093.000000000,-184.91
1094.000000000,-184.44
1095.000000000,-184.17
1096.000000000,-184.01
1097.000000000,-183.97
1098.000000000,-184.59
1099.000000000,-184.10
1100.000000000,-183.96
1101.000000000,-183.87
1102.000000000,-183.82
1103.000000000,-183.79
1104.000000000,-183.76
1105.000000000,-183.75
1106.000000000,-183.74
1107.000000000,-183.73
1108.000000000,-183.72
1109.000000000,-183.71
1110.000000000,-183.71
1111.000000000,-183.70
1112.000000000,-183.70
1113.000000000,-183.70
1114.000000000,-183.69
1115.000000000,-183.69
1116.000000000,-183.68
1117.000000000,-183.68
1118.000000000,-183.67
1119.000000000,-183.67
1120.000000000,-183.66
1121.000000000,-183.66
1122.000000000,-186.05
1123.000000000,-184.57
1124.000000000,-184.18
1125.000000000,-183.97
1126.000000000,-183.85
1127.000000000,-183.77
1128.000000000,-183.72
1129.000000000,-183.69
1130.000000000,-183.67
1131.000000000,-183.65
1132.000000000,-183.64
1133.000000000,-183.64
1134.000000000,-183.63
1135.000000000,-183.62
1136.000000000,-183.62
1137.000000000,-183.61
1138.000000000,-183.61
1139.000000000,-183.61
1140.000000000,-183.60
1141.000000000,-183.60
1142.000000000,-183.59
1143.000000000,-183.59
1144.000000000,-183.59
1145.000000000,-183.58
1146.000000000,-183.58
1147.000000000,-183.58
1148.000000000,-184.49
1149.000000000,-186.45
1150.000000000,-184.75
1151.000000000,-184.25
1152.000000000,-183.99
1153.000000000,-183.83
1154.000000000,-183.73
1155.000000000,-183.68
1156.000000000,-183.64
1157.000000000,-183.61
1158.000000000,-183.59
1159.000000000,-183.58
1160.000000000,-183.57
1161.000000000,-183.56
1162.000000000,-183.55
1163.000000000,-187.77
1164.000000000,-187.85
1165.000000000,-189.51
1166.000000000,-190.22
1167.000000000,-189.12
1168.000000000,-186.38
1169.000000000,-185.29
1170.000000000,-184.67
1171.000000000,-184.29
1172.000000000,-184.14
1173.000000000,-183.94
1174.000000000,-185.79
1175.000000000,-184.52
1176.000000000,-184.15
1177.000000000,-183.95
1178.000000000,-183.83
1179.000000000,-184.01
1180.000000000,-183.80
1181.000000000,-183.73
1182.000000000,-183.68
1183.000000000,-183.65
1184.000000000,-183.63
1185.000000000,-183.61
1186.000000000,-183.60
1187.000000000,-183.63
1188.000000000,-183.60
1189.000000000,-183.59
1190.000000000,-183.58
1191.000000000,-183.57
1192.000000000,-183.56
1193.000000000,-183.55
1194.000000000,-183.55
1195.000000000,-183.54
1196.000000000,-183.54
1197.000000000,-183.60
1198.000000000,-183.55
1199.000000000,-185.28
1200.000000000,-184.20
1201.000000000,-183.91
1202.000000000,-183.75
1203.000000000,-195.22
1204.000000000,-190.61
1205.000000000,-187.20
1206.000000000,-185.79
1207.000000000,-184.95
1208.000000000,-184.49
1209.000000000,-184.16
1210.000000000,-184.14
1211.000000000,-183.91
1212.000000000,-183.79
1213.000000000,-184.87
1214.000000000,-184.11
1215.000000000,-183.89
1216.000000000,-183.80
1217.000000000,-183.71
1218.000000000,-183.70
1219.000000000,-183.64
1220.000000000,-183.61
1221.000000000,-183.59
1222.000000000,-183.57
1223.000000000,-183.56
1224.000000000,-183.55
1225.000000000,-183.92
1226.000000000,-183.68
1227.000000000,-183.61
1228.000000000,-183.57
1229.000000000,-183.60
1230.000000000,-183.56
1231.000000000,-184.14
1232.000000000,-184.13
1233.000000000,-183.81
1234.000000000,-185.08
1235.000000000,-187.82
1236.000000000,-186.03
1237.000000000,-184.84
1238.000000000,-184.32
1239.000000000,-184.02
1240.000000000,-183.84
1241.000000000,-183.73
1242.000000000,-183.66
1243.000000000,-183.64
1244.000000000,-183.59
1245.000000000,-183.56
1246.000000000,-183.71
1247.000000000,-183.60
1248.000000000,-183.98
1249.000000000,-191.21
1250.000000000,-188.16
1251.000000000,-186.04
1252.000000000,-185.00
1253.000000000,-184.45
1254.000000000,-184.12
1255.000000000,-183.92
1256.000000000,-183.79
1257.000000000,-183.71
1258.000000000,-183.65
1259.000000000,-183.62
1260.000000000,-183.67
1261.000000000,-183.60
1262.000000000,-183.58
1263.000000000,-183.56
1264.000000000,-183.55
1265.000000000,-183.54
1266.000000000,-183.53
1267.000000000,-185.19
1268.000000000,-184.16
1269.000000000,-183.88
1270.000000000,-183.74
1271.000000000,-183.65
1272.000000000,-183.59
1273.000000000,-185.17
1274.000000000,-196.72
1275.000000000,-189.18
1276.000000000,-186.86
1277.000000000,-185.53
1278.000000000,-184.80
1279.000000000,-184.36
1280.000000000,-184.09
1281.000000000,-183.92
1282.000000000,-183.81
1283.000000000,-183.73
1284.000000000,-183.68
1285.000000000,-183.65
1286.000000000,-183.62
1287.000000000,-183.62
1288.000000000,-183.60
1289.000000000,-183.58
1290.000000000,-183.57
1291.000000000,-183.56
1292.000000000,-183.56
1293.000000000,-183.55
1294.000000000,-183.55
1295.000000000,-183.54
1296.000000000,-183.54
1297.000000000,-183.53
1298.000000000,-183.53
1299.000000000,-183.52
1300.000000000,-183.52
1301.000000000,-183.52
1302.000000000,-183.51
1303.000000000,-183.55
1304.000000000,-184.83
1305.000000000,-184.14
1306.000000000,-183.85
1307.000000000,-183.77
1308.000000000,-183.65
1309.000000000,-183.59
1310.000000000,-183.56
1311.000000000,-183.53
1312.000000000,-183.51
1313.000000000,-183.50
1314.000000000,-183.49
1315.000000000,-183.48
1316.000000000,-183.48
1317.000000000,-183.47
1318.000000000,-183.47
1319.000000000,-183.46
1320.000000000,-183.46
1321.000000000,-188.06
1322.000000000,-189.21
1323.000000000,-187.53
1324.000000000,-185.86
1325.000000000,-187.66
1326.000000000,-186.29
1327.000000000,-185.33
1328.000000000,-194.25
1329.000000000,-189.13
1330.000000000,-188.45
1331.000000000,-188.42
1332.000000000,-186.03
1333.000000000,-185.40
1334.000000000,-184.67
1335.000000000,-184.29
1336.000000000,-184.22
1337.000000000,-184.68
1338.000000000,-184.44
1339.000000000,-184.71
1340.000000000,-184.53
1341.000000000,-184.48
1342.000000000,-185.46
1343.000000000,-184.45
1344.000000000,-184.11
1345.000000000,-183.93
1346.000000000,-183.81
1347.000000000,-183.74
1348.000000000,-183.69
1349.000000000,-183.66
1350.000000000,-184.13
1351.000000000,-183.81
1352.000000000,-184.99
1353.000000000,-184.28
1354.000000000,-184.53
1355.000000000,-184.03
1356.000000000,-183.85
1357.000000000,-183.75
1358.000000000,-183.69
1359.000000000,-183.65
1360.000000000,-183.62
1361.000000000,-183.60
1362.000000000,-183.58
1363.000000000,-183.57
1364.000000000,-189.65
1365.000000000,-199.89
1366.000000000,-191.84
1367.000000000,-188.10
1368.000000000,-186.34
1369.000000000,-185.34
1370.000000000,-184.74
1371.000000000,-184.37
1372.000000000,-184.14
1373.000000000,-183.99
1374.000000000,-183.89
1375.000000000,-183.82
1376.000000000,-183.77
1377.000000000,-183.77
1378.000000000,-183.72
1379.000000000,-183.70
1380.000000000,-183.68
1381.000000000,-183.66
1382.000000000,-183.65
1383.000000000,-183.64
1384.000000000,-183.63
1385.000000000,-183.63
1386.000000000,-183.62
1387.000000000,-183.61
1388.000000000,-183.61
1389.000000000,-183.60
1390.000000000,-183.62
1391.000000000,-183.60
1392.000000000,-183.59
1393.000000000,-183.58
1394.000000000,-183.57
1395.000000000,-183.57
1396.000000000,-183.56
1397.000000000,-183.55
1398.000000000,-183.55
1399.000000000,-183.54
1400.000000000,-183.54
1401.000000000,-183.53
1402.000000000,-183.53
1403.000000000,-183.52
1404.000000000,-186.19
1405.000000000,-184.64
1406.000000000,-184.19
1407.000000000,-184.27
1408.000000000,-183.90
1409.000000000,-183.75
1410.000000000,-187.67
1411.000000000,-185.27
1412.000000000,-184.51
1413.000000000,-184.12
1414.000000000,-183.89
1415.000000000,-183.75
1416.000000000,-183.66
1417.000000000,-183.61
1418.000000000,-183.57
1419.000000000,-183.54
1420.000000000,-183.52
1421.000000000,-183.50
1422.000000000,-183.49
1423.000000000,-183.48
1424.000000000,-183.47
1425.000000000,-183.47
1426.000000000,-183.82
1427.000000000,-183.60
1428.000000000,-183.53
1429.000000000,-183.49
1430.000000000,-183.47
1431.000000000,-183.45
1432.000000000,-183.44
1433.000000000,-184.97
1434.000000000,-186.62
1435.000000000,-193.50
1436.000000000,-188.44
1437.000000000,-186.19
1438.000000000,-185.12
1439.000000000,-184.51
1440.000000000,-184.14
1441.000000000,-183.92
1442.000000000,-183.77
1443.000000000,-183.89
1444.000000000,-183.70
1445.000000000,-183.62
1446.000000000,-183.61
1447.000000000,-183.56
1448.000000000,-183.53
1449.000000000,-183.51
1450.000000000,-183.49
1451.000000000,-183.48
1452.000000000,-183.68
1453.000000000,-183.55
1454.000000000,-183.87
1455.000000000,-183.63
1456.000000000,-183.55
1457.000000000,-183.51
1458.000000000,-183.48
1459.000000000,-183.47
1460.000000000,-183.54
1461.000000000,-183.50
1462.000000000,-183.47
1463.000000000,-183.67
1464.000000000,-183.53
1465.000000000,-183.48
1466.000000000,-183.46
1467.000000000,-183.44
1468.000000000,-183.43
1469.000000000,-183.42
1470.000000000,-183.42
1471.000000000,-183.41
1472.000000000,-183.41
1473.000000000,-183.40
1474.000000000,-183.40
1475.000000000,-183.73
1476.000000000,-184.18
1477.000000000,-185.16
1478.000000000,-184.14
1479.000000000,-185.67
1480.000000000,-184.37
1481.000000000,-183.97
1482.000000000,-183.75
1483.000000000,-183.62
1484.000000000,-183.54
1485.000000000,-183.49
1486.000000000,-183.46
1487.000000000,-183.44
1488.000000000,-183.42
1489.000000000,-183.52
1490.000000000,-183.45
1491.000000000,-183.42
1492.000000000,-183.41
1493.000000000,-183.40
1494.000000000,-183.39
1495.000000000,-183.39
1496.000000000,-183.38
1497.000000000,-183.44
1498.000000000,-183.40
1499.000000000,-183.39
1500.000000000,-183.38
1501.000000000,-183.37
1502.000000000,-183.37
1503.000000000,-183.36
1504.000000000,-183.36
1505.000000000,-183.36
1506.000000000,-189.28
1507.000000000,-185.63
1508.000000000,-184.67
1509.000000000,-184.27
1510.000000000,-183.90
1511.000000000,-183.71
1512.000000000,-184.38
1513.000000000,-183.82
1514.000000000,-183.65
1515.000000000,-183.55
1516.000000000,-183.48
1517.000000000,-183.44
1518.000000000,-183.42
1519.000000000,-183.40
1520.000000000,-183.39
1521.000000000,-183.38
1522.000000000,-183.37
1523.000000000,-183.36
1524.000000000,-183.36
1525.000000000,-183.76
1526.000000000,-183.51
1527.000000000,-183.44
1528.000000000,-183.40
1529.000000000,-183.38
1530.000000000,-183.36
1531.000000000,-183.45
1532.000000000,-183.39
1533.000000000,-183.36
1534.000000000,-183.35
1535.000000000,-183.34
1536.000000000,-183.33
1537.000000000,-183.33
1538.000000000,-183.32
1539.000000000,-183.32
1540.000000000,-183.31
1541.000000000,-183.31
1542.000000000,-183.30
1543.000000000,-183.30
1544.000000000,-183.37
1545.000000000,-183.32
1546.000000000,-183.30
1547.000000000,-183.29
1548.000000000,-183.28
1549.000000000,-185.91
1550.000000000,-184.29
1551.000000000,-183.85
1552.000000000,-183.62
1553.000000000,-188.49
1554.000000000,-185.33
1555.000000000,-184.47
1556.000000000,-184.01
1557.000000000,-183.74
1558.000000000,-183.57
1559.000000000,-183.47
1560.000000000,-183.40
1561.000000000,-183.36
1562.000000000,-184.96
1563.000000000,-184.39
1564.000000000,-184.36
1565.000000000,-186.05
1566.000000000,-184.46
1567.000000000,-184.13
1568.000000000,-184.53
1569.000000000,-183.88
1570.000000000,-183.64
1571.000000000,-183.51
1572.000000000,-183.42
1573.000000000,-183.37
1574.000000000,-183.33
1575.000000000,-183.31
1576.000000000,-183.29
1577.000000000,-183.27
1578.000000000,-183.26
1579.000000000,-183.25
1580.000000000,-183.25
1581.000000000,-183.24
1582.000000000,-183.23
1583.000000000,-183.23
1584.000000000,-183.22
1585.000000000,-183.22
1586.000000000,-183.22
1587.000000000,-183.21
1588.000000000,-183.21
1589.000000000,-183.20
1590.000000000,-183.20
1591.000000000,-183.19
1592.000000000,-185.27
1593.000000000,-183.99
1594.000000000,-183.65
1595.000000000,-183.46
1596.000000000,-183.36
1597.000000000,-183.29
1598.000000000,-183.30
1599.000000000,-183.24
1600.000000000,-183.22
1601.000000000,-187.26
1602.000000000,-185.02
1603.000000000,-187.54
1604.000000000,-185.12
1605.000000000,-184.44
1606.000000000,-183.94
1607.000000000,-183.66
1608.000000000,-183.50
1609.000000000,-183.39
1610.000000000,-187.41
1611.000000000,-184.93
1612.000000000,-197.52
1613.000000000,-190.49
1614.000000000,-187.48
1615.000000000,-186.67
1616.000000000,-187.48
1617.000000000,-185.67
1618.000000000,-184.69
1619.000000000,-184.19
1620.000000000,-183.88
1621.000000000,-183.69
1622.000000000,-183.57
1623.000000000,-183.49
1624.000000000,-183.43
1625.000000000,-183.39
1626.000000000,-183.37
1627.000000000,-183.35
1628.000000000,-183.35
1629.000000000,-183.32
1630.000000000,-183.31
1631.000000000,-183.30
1632.000000000,-183.29
1633.000000000,-183.29
1634.000000000,-183.28
1635.000000000,-183.27
1636.000000000,-183.32
1637.000000000,-183.29
1638.000000000,-183.30
1639.000000000,-184.40
1640.000000000,-183.92
1641.000000000,-183.59
1642.000000000,-183.45
1643.000000000,-183.37
1644.000000000,-183.33
1645.000000000,-183.29
1646.000000000,-183.27
1647.000000000,-183.39
1648.000000000,-183.47
1649.000000000,-184.89
1650.000000000,-185.84
1651.000000000,-184.36
1652.000000000,-183.89
1653.000000000,-183.63
1654.000000000,-183.48
1655.000000000,-183.41
1656.000000000,-183.66
1657.000000000,-184.13
1658.000000000,-184.72
1659.000000000,-184.40
1660.000000000,-184.05
1661.000000000,-183.86
1662.000000000,-183.57
1663.000000000,-183.43
1664.000000000,-183.35
1665.000000000,-183.31
1666.000000000,-187.16
1667.000000000,-184.77
1668.000000000,-184.10
1669.000000000,-183.75
1670.000000000,-183.55
1671.000000000,-183.42
1672.000000000,-183.35
1673.000000000,-183.76
1674.000000000,-183.67
1675.000000000,-184.10
1676.000000000,-184.36
1677.000000000,-183.73
1678.000000000,-183.58
1679.000000000,-183.42
1680.000000000,-183.33
1681.000000000,-183.52
1682.000000000,-188.35
1683.000000000,-185.21
1684.000000000,-184.41
1685.000000000,-183.92
1686.000000000,-183.65
1687.000000000,-183.49
1688.000000000,-183.38
1689.000000000,-183.68
1690.000000000,-183.59
1691.000000000,-183.39
1692.000000000,-183.32
1693.000000000,-183.27
1694.000000000,-183.23
1695.000000000,-183.21
1696.000000000,-183.19
1697.000000000,-184.41
1698.000000000,-185.15
1699.000000000,-184.20
1700.000000000,-184.68
1701.000000000,-183.88
1702.000000000,-183.59
1703.000000000,-183.42
1704.000000000,-183.32
1705.000000000,-183.26
1706.000000000,-183.22
1707.000000000,-183.19
1708.000000000,-183.23
1709.000000000,-183.18
1710.000000000,-183.18
1711.000000000,-183.15
1712.000000000,-183.14
1713.000000000,-183.12
1714.000000000,-183.11
1715.000000000,-183.11
1716.000000000,-183.10
1717.000000000,-183.09
1718.000000000,-183.09
1719.000000000,-183.08
1720.000000000,-183.08
1721.000000000,-183.07
1722.000000000,-183.07
1723.000000000,-183.06
1724.000000000,-183.15
1725.000000000,-183.09
1726.000000000,-183.08
1727.000000000,-183.14
1728.000000000,-183.08
1729.000000000,-187.44
1730.000000000,-187.32
1731.000000000,-193.81
1732.000000000,-196.27
1733.000000000,-192.98
1734.000000000,-189.38
1735.000000000,-187.08
1736.000000000,-185.50
1737.000000000,-184.66
1738.000000000,-186.71
1739.000000000,-185.24
1740.000000000,-184.36
1741.000000000,-183.94
1742.000000000,-183.69
1743.000000000,-183.53
1744.000000000,-184.78
1745.000000000,-183.96
1746.000000000,-183.65
1747.000000000,-183.49
1748.000000000,-183.39
1749.000000000,-183.33
1750.000000000,-183.31
1751.000000000,-183.27
1752.000000000,-183.24
1753.000000000,-183.23
1754.000000000,-183.21
1755.000000000,-183.20
1756.000000000,-183.19
1757.000000000,-183.19
1758.000000000,-183.18
1759.000000000,-183.17
1760.000000000,-183.17
1761.000000000,-183.16
1762.000000000,-183.16
1763.000000000,-183.15
1764.000000000,-183.15
1765.000000000,-183.14
1766.000000000,-183.16
1767.000000000,-183.14
1768.000000000,-183.14
1769.000000000,-183.13
1770.000000000,-183.12
1771.000000000,-183.12
1772.000000000,-183.12
1773.000000000,-183.11
1774.000000000,-183.16
1775.000000000,-183.13
1776.000000000,-183.12
1777.000000000,-183.51
1778.000000000,-183.26
1779.000000000,-183.30
1780.000000000,-183.20
1781.000000000,-183.15
1782.000000000,-183.13
1783.000000000,-183.11
1784.000000000,-183.10
1785.000000000,-183.09
1786.000000000,-183.08
1787.000000000,-183.07
1788.000000000,-183.07
1789.000000000,-183.06
1790.000000000,-183.06
1791.000000000,-183.06
1792.000000000,-183.05
1793.000000000,-183.05
1794.000000000,-183.05
1795.000000000,-183.04
1796.000000000,-183.04
1797.000000000,-183.03
1798.000000000,-183.03
1799.000000000,-183.03
1800.000000000,-183.02
1801.000000000,-184.20
1802.000000000,-187.77
1803.000000000,-186.13
1804.000000000,-184.59
1805.000000000,-183.97
1806.000000000,-183.62
1807.000000000,-183.41
1808.000000000,-183.28
1809.000000000,-183.19
1810.000000000,-183.14
1811.000000000,-183.27
1812.000000000,-184.67
1813.000000000,-183.69
1814.000000000,-183.73
1815.000000000,-183.40
1816.000000000,-183.25
1817.000000000,-183.17
1818.000000000,-183.16
1819.000000000,-183.10
1820.000000000,-183.07
1821.000000000,-183.05
1822.000000000,-183.20
1823.000000000,-183.18
1824.000000000,-183.09
1825.000000000,-183.08
1826.000000000,-183.04
1827.000000000,-183.02
1828.000000000,-183.06
1829.000000000,-183.02
1830.000000000,-183.01
1831.000000000,-183.00
1832.000000000,-182.99
1833.000000000,-182.98
1834.000000000,-182.98
1835.000000000,-182.97
1836.000000000,-182.97
1837.000000000,-182.96
1838.000000000,-182.96
1839.000000000,-182.96
1840.000000000,-182.95
1841.000000000,-182.95
1842.000000000,-183.03
1843.000000000,-182.98
1844.000000000,-182.96
1845.000000000,-183.02
1846.000000000,-183.02
1847.000000000,-182.97
1848.000000000,-182.95
1849.000000000,-182.94
1850.000000000,-182.93
1851.000000000,-182.93
1852.000000000,-182.92
1853.000000000,-182.91
1854.000000000,-182.91
1855.000000000,-182.91
1856.000000000,-182.90
1857.000000000,-182.90
1858.000000000,-182.89
1859.000000000,-182.89
1860.000000000,-182.98
1861.000000000,-182.92
1862.000000000,-182.90
1863.000000000,-182.89
1864.000000000,-182.93
1865.000000000,-182.90
1866.000000000,-182.88
1867.000000000,-182.87
1868.000000000,-182.87
1869.000000000,-182.86
1870.000000000,-183.15
1871.000000000,-183.06
1872.000000000,-182.95
1873.000000000,-182.90
1874.000000000,-182.87
1875.000000000,-182.86
1876.000000000,-183.27
1877.000000000,-184.24
1878.000000000,-188.38
1879.000000000,-185.43
1880.000000000,-184.29
1881.000000000,-183.82
1882.000000000,-183.43
1883.000000000,-183.21
1884.000000000,-183.08
1885.000000000,-183.00
1886.000000000,-183.20
1887.000000000,-183.01
1888.000000000,-182.94
1889.000000000,-182.90
1890.000000000,-182.88
1891.000000000,-182.86
1892.000000000,-182.85
1893.000000000,-182.84
1894.000000000,-182.83
1895.000000000,-182.83
1896.000000000,-182.82
1897.000000000,-182.82
1898.000000000,-182.82
1899.000000000,-182.81
1900.000000000,-182.81
1901.000000000,-182.81
1902.000000000,-182.81
1903.000000000,-182.80
1904.000000000,-182.80
1905.000000000,-182.80
1906.000000000,-182.80
1907.000000000,-182.79
1908.000000000,-182.79
1909.000000000,-182.79
1910.000000000,-182.78
1911.000000000,-182.78
1912.000000000,-182.78
1913.000000000,-183.02
1914.000000000,-182.87
1915.000000000,-182.83
1916.000000000,-182.80
1917.000000000,-182.78
1918.000000000,-182.77
1919.000000000,-182.77
1920.000000000,-182.76
1921.000000000,-182.75
1922.000000000,-182.75
1923.000000000,-182.74
1924.000000000,-182.74
1925.000000000,-182.74
1926.000000000,-182.73
1927.000000000,-182.73
1928.000000000,-182.73
1929.000000000,-182.72
1930.000000000,-182.85
1931.000000000,-182.77
1932.000000000,-182.75
1933.000000000,-182.73
1934.000000000,-182.72
1935.000000000,-182.71
1936.000000000,-182.71
1937.000000000,-182.72
1938.000000000,-182.79
1939.000000000,-182.73
1940.000000000,-182.71
1941.000000000,-182.70
1942.000000000,-183.51
1943.000000000,-183.00
1944.000000000,-182.86
1945.000000000,-182.79
1946.000000000,-182.74
1947.000000000,-182.72
1948.000000000,-182.70
1949.000000000,-182.94
1950.000000000,-188.48
1951.000000000,-185.82
1952.000000000,-184.32
1953.000000000,-183.66
1954.000000000,-183.29
1955.000000000,-183.07
1956.000000000,-182.94
1957.000000000,-182.85
1958.000000000,-182.79
1959.000000000,-182.76
1960.000000000,-182.73
1961.000000000,-182.71
1962.000000000,-182.70
1963.000000000,-182.69
1964.000000000,-182.72
1965.000000000,-182.69
1966.000000000,-183.21
1967.000000000,-188.35
1968.000000000,-185.02
1969.000000000,-184.00
1970.000000000,-183.48
1971.000000000,-183.18
1972.000000000,-183.00
1973.000000000,-182.88
1974.000000000,-182.81
1975.000000000,-182.76
1976.000000000,-182.73
1977.000000000,-182.71
1978.000000000,-182.69
1979.000000000,-182.68
1980.000000000,-182.67
1981.000000000,-182.95
1982.000000000,-182.77
1983.000000000,-182.72
1984.000000000,-182.69
1985.000000000,-182.67
1986.000000000,-182.65
1987.000000000,-182.64
1988.000000000,-182.65
1989.000000000,-182.64
1990.000000000,-182.63
1991.000000000,-182.62
1992.000000000,-182.62
1993.000000000,-182.61
1994.000000000,-182.61
1995.000000000,-182.63
1996.000000000,-182.99
1997.000000000,-182.75
1998.000000000,-182.69
1999.000000000,-182.72
2000.000000000,-182.66
2001.000000000,-182.63
2002.000000000,-182.61
2003.000000000,-182.60
2004.000000000,-182.60
2005.000000000,-182.58
2006.000000000,-182.58
2007.000000000,-182.89
2008.000000000,-182.69
2009.000000000,-182.64
2010.000000000,-182.61
2011.000000000,-182.59
2012.000000000,-183.15
2013.000000000,-183.79
2014.000000000,-185.41
2015.000000000,-186.22
2016.000000000,-185.25
2017.000000000,-185.67
2018.000000000,-184.07
2019.000000000,-183.48
2020.000000000,-183.14
2021.000000000,-182.94
2022.000000000,-182.81
2023.000000000,-182.73
2024.000000000,-182.68
2025.000000000,-182.64
2026.000000000,-182.62
2027.000000000,-182.60
2028.000000000,-182.58
2029.000000000,-182.57
2030.000000000,-182.56
2031.000000000,-182.56
2032.000000000,-182.55
2033.000000000,-182.54
2034.000000000,-182.54
2035.000000000,-182.53
2036.000000000,-182.53
2037.000000000,-182.53
2038.000000000,-188.14
2039.000000000,-184.84
2040.000000000,-183.83
2041.000000000,-183.32
2042.000000000,-183.02
2043.000000000,-182.84
2044.000000000,-182.73
2045.000000000,-182.66
2046.000000000,-182.62
2047.000000000,-182.59
2048.000000000,-182.59
2049.000000000,-184.69
2050.000000000,-184.85
2051.000000000,-185.55
2052.000000000,-184.38
2053.000000000,-183.53
2054.000000000,-183.14
2055.000000000,-182.92
2056.000000000,-182.78
2057.000000000,-182.69
2058.000000000,-183.10
2059.000000000,-183.68
2060.000000000,-183.03
2061.000000000,-182.82
2062.000000000,-182.71
2063.000000000,-182.64
2064.000000000,-182.59
2065.000000000,-182.56
2066.000000000,-182.54
2067.000000000,-182.53
2068.000000000,-182.52
2069.000000000,-182.51
