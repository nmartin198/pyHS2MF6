time,FINEGAN,704,703,DOLAN,701
1.000000000000,-0.11361E+06,-0.12836E+06,-84869.,-14619.,-16610.
2.000000000000,-0.12433E+06,-0.12737E+06,-78981.,-14626.,-16628.
3.000000000000,-0.12269E+06,-0.12107E+06,-71976.,-14631.,-16640.
4.000000000000,-0.11862E+06,-0.11501E+06,-66338.,-14636.,-16650.
5.000000000000,-0.11426E+06,-0.10957E+06,-61696.,-14640.,-16659.
6.000000000000,-0.11010E+06,-0.10470E+06,-57727.,-14643.,-16664.
7.000000000000,-0.10623E+06,-0.10032E+06,-54248.,-14646.,-16668.
8.000000000000,-0.10263E+06,-96332.,-51144.,-14647.,-16671.
9.000000000000,-99311.,-92694.,-48356.,-14649.,-16673.
10.00000000000,-96221.,-89342.,-45823.,-14649.,-16675.
11.00000000000,-93318.,-86222.,-43492.,-14650.,-16677.
12.00000000000,-90594.,-83320.,-41350.,-14650.,-16678.
13.00000000000,-88037.,-80610.,-39377.,-14650.,-16678.
14.00000000000,-85632.,-78073.,-37554.,-14650.,-16678.
15.00000000000,-83365.,-75690.,-35864.,-14650.,-16678.
16.00000000000,-81225.,-73447.,-34296.,-14650.,-16677.
17.00000000000,-79199.,-71332.,-32836.,-14650.,-16677.
18.00000000000,-77280.,-69332.,-31475.,-14650.,-16677.
19.00000000000,-75458.,-67439.,-30204.,-14650.,-16677.
20.00000000000,-73727.,-65644.,-29016.,-14650.,-16676.
21.00000000000,-72078.,-63939.,-27902.,-14650.,-16676.
22.00000000000,-70507.,-62318.,-26859.,-14650.,-16675.
23.00000000000,-69008.,-60775.,-25878.,-14649.,-16675.
24.00000000000,-67574.,-59303.,-24956.,-14649.,-16674.
25.00000000000,-66203.,-57899.,-24089.,-14649.,-16674.
26.00000000000,-64889.,-56557.,-23271.,-14648.,-16673.
27.00000000000,-63629.,-55273.,-22499.,-14648.,-16672.
28.00000000000,-62419.,-54044.,-21770.,-14647.,-16672.
29.00000000000,-61256.,-52866.,-21081.,-14647.,-16671.
30.00000000000,-60137.,-51736.,-20429.,-14647.,-16670.
31.00000000000,-59060.,-50651.,-19811.,-14646.,-16670.
32.00000000000,-58021.,-49609.,-19225.,-14646.,-16669.
33.00000000000,-57018.,-48607.,-18669.,-14645.,-16668.
34.00000000000,-56050.,-47642.,-18140.,-14645.,-16668.
35.00000000000,-55114.,-46713.,-17638.,-14644.,-16667.
36.00000000000,-54209.,-45818.,-17160.,-14644.,-16666.
37.00000000000,-53333.,-44954.,-16705.,-14644.,-16666.
38.00000000000,-52484.,-44121.,-16271.,-14643.,-16665.
39.00000000000,-51661.,-43317.,-15857.,-14643.,-16665.
40.00000000000,-50862.,-42539.,-15461.,-14642.,-16664.
41.00000000000,-50087.,-41788.,-15084.,-14642.,-16663.
42.00000000000,-49335.,-41061.,-14723.,-14642.,-16663.
43.00000000000,-48603.,-40357.,-14378.,-14641.,-16662.
44.00000000000,-47892.,-39676.,-14047.,-14641.,-16662.
45.00000000000,-47200.,-39015.,-13730.,-14640.,-16661.
46.00000000000,-46526.,-38376.,-13427.,-14640.,-16661.
47.00000000000,-45870.,-37755.,-13136.,-14640.,-16660.
48.00000000000,-45231.,-37153.,-12856.,-14639.,-16660.
49.00000000000,-44607.,-36569.,-12588.,-14639.,-16659.
50.00000000000,-44000.,-36002.,-12330.,-14639.,-16659.
51.00000000000,-43407.,-35450.,-12082.,-14638.,-16658.
52.00000000000,-42829.,-34916.,-11843.,-14638.,-16658.
53.00000000000,-42264.,-34395.,-11614.,-14638.,-16657.
54.00000000000,-41712.,-33889.,-11392.,-14637.,-16657.
55.00000000000,-41173.,-33396.,-11179.,-14637.,-16656.
56.00000000000,-40647.,-32917.,-10974.,-14637.,-16656.
57.00000000000,-40132.,-32450.,-10776.,-14636.,-16655.
58.00000000000,-39628.,-31996.,-10584.,-14636.,-16655.
59.00000000000,-39136.,-31553.,-10400.,-14636.,-16654.
60.00000000000,-38654.,-31121.,-10221.,-14635.,-16654.
61.00000000000,-38182.,-30700.,-10049.,-14635.,-16653.
62.00000000000,-37720.,-30290.,-9881.8,-14635.,-16653.
63.00000000000,-37267.,-29890.,-9720.5,-14634.,-16652.
64.00000000000,-36824.,-29500.,-9564.5,-14634.,-16652.
65.00000000000,-36391.,-29118.,-9413.4,-14634.,-16652.
66.00000000000,-35965.,-28746.,-9267.1,-14634.,-16651.
67.00000000000,-35549.,-28383.,-9125.3,-14633.,-16651.
68.00000000000,-35140.,-28028.,-8987.9,-14633.,-16650.
69.00000000000,-34741.,-27683.,-8856.0,-14633.,-16650.
70.00000000000,-34349.,-27344.,-8726.6,-14632.,-16650.
71.00000000000,-33964.,-27013.,-8601.1,-14632.,-16649.
72.00000000000,-33586.,-26689.,-8479.2,-14632.,-16649.
73.00000000000,-33215.,-26373.,-8360.9,-14632.,-16648.
74.00000000000,-32852.,-26063.,-8246.0,-14631.,-16648.
75.00000000000,-32495.,-25760.,-8134.4,-14631.,-16648.
76.00000000000,-32144.,-25464.,-8026.0,-14631.,-16647.
77.00000000000,-31800.,-25173.,-7920.5,-14631.,-16647.
78.00000000000,-31463.,-24889.,-7818.0,-14630.,-16647.
79.00000000000,-31131.,-24611.,-7718.2,-14630.,-16646.
80.00000000000,-30805.,-24339.,-7621.1,-14630.,-16646.
81.00000000000,-30486.,-24072.,-7526.6,-14630.,-16645.
82.00000000000,-30172.,-23812.,-7435.3,-14629.,-16645.
83.00000000000,-29864.,-23556.,-7345.6,-14629.,-16645.
84.00000000000,-29561.,-23305.,-7258.1,-14629.,-16644.
85.00000000000,-29263.,-23059.,-7172.9,-14629.,-16644.
86.00000000000,-28971.,-22818.,-7089.9,-14629.,-16644.
87.00000000000,-28683.,-22582.,-7008.9,-14628.,-16643.
88.00000000000,-28400.,-22350.,-6930.0,-14628.,-16643.
89.00000000000,-28122.,-22123.,-6853.0,-14628.,-16642.
90.00000000000,-27849.,-21900.,-6777.8,-14628.,-16642.
91.00000000000,-27581.,-21681.,-6704.5,-14628.,-16641.
92.00000000000,-27317.,-21467.,-6632.8,-14628.,-16641.
93.00000000000,-27061.,-21260.,-6565.7,-14627.,-16640.
94.00000000000,-26807.,-21053.,-6497.3,-14627.,-16640.
95.00000000000,-26556.,-20850.,-6430.1,-14627.,-16639.
96.00000000000,-26309.,-20650.,-6364.6,-14627.,-16639.
97.00000000000,-26066.,-20455.,-6300.6,-14627.,-16638.
98.00000000000,-25826.,-20262.,-6238.0,-14627.,-16638.
99.00000000000,-25591.,-20074.,-6177.0,-14626.,-16637.
100.0000000000,-25360.,-19889.,-6117.2,-14626.,-16637.
101.0000000000,-25132.,-19707.,-6058.9,-14626.,-16636.
102.0000000000,-24908.,-19528.,-6001.7,-14626.,-16636.
103.0000000000,-24687.,-19352.,-5945.8,-14626.,-16635.
104.0000000000,-24470.,-19179.,-5891.2,-14626.,-16635.
105.0000000000,-24256.,-19010.,-5837.6,-14625.,-16635.
106.0000000000,-24046.,-18843.,-5785.2,-14625.,-16634.
107.0000000000,-23839.,-18679.,-5733.9,-14625.,-16634.
108.0000000000,-23637.,-18520.,-5685.1,-14625.,-16633.
109.0000000000,-23437.,-18362.,-5635.8,-14625.,-16633.
110.0000000000,-23240.,-18206.,-5587.3,-14625.,-16632.
111.0000000000,-23045.,-18052.,-5539.8,-14624.,-16632.
112.0000000000,-22853.,-17901.,-5493.4,-14624.,-16631.
113.0000000000,-22664.,-17753.,-5447.8,-14624.,-16631.
114.0000000000,-22478.,-17607.,-5403.2,-14624.,-16631.
115.0000000000,-22295.,-17464.,-5359.4,-14624.,-16630.
116.0000000000,-22115.,-17323.,-5316.5,-14624.,-16630.
117.0000000000,-21937.,-17184.,-5274.5,-14624.,-16629.
118.0000000000,-21769.,-17054.,-5238.0,-14623.,-16629.
119.0000000000,-21612.,-16931.,-5205.4,-14623.,-16628.
120.0000000000,-21445.,-16796.,-5164.5,-14623.,-16628.
121.0000000000,-21278.,-16664.,-5123.8,-14623.,-16628.
122.0000000000,-21117.,-16538.,-5087.1,-14623.,-16627.
123.0000000000,-20955.,-16411.,-5048.3,-14623.,-16627.
124.0000000000,-20794.,-16285.,-5010.1,-14623.,-16626.
125.0000000000,-20636.,-16161.,-4972.9,-14623.,-16626.
126.0000000000,-20479.,-16040.,-4936.5,-14622.,-16626.
127.0000000000,-20325.,-15921.,-4900.9,-14622.,-16625.
128.0000000000,-20173.,-15803.,-4866.0,-14622.,-16625.
129.0000000000,-20024.,-15688.,-4831.9,-14622.,-16624.
130.0000000000,-19879.,-15576.,-4799.8,-14622.,-16624.
131.0000000000,-19737.,-15467.,-4768.7,-14622.,-16623.
132.0000000000,-19594.,-15356.,-4736.1,-14622.,-16623.
133.0000000000,-19453.,-15246.,-4703.9,-14621.,-16623.
134.0000000000,-19314.,-15139.,-4672.4,-14621.,-16622.
135.0000000000,-19180.,-15037.,-4643.9,-14621.,-16622.
136.0000000000,-19045.,-14932.,-4613.5,-14621.,-16621.
137.0000000000,-18912.,-14829.,-4583.4,-14621.,-16621.
138.0000000000,-18780.,-14727.,-4553.9,-14621.,-16621.
139.0000000000,-18650.,-14628.,-4525.0,-14621.,-16620.
140.0000000000,-18521.,-14529.,-4496.6,-14620.,-16620.
141.0000000000,-18395.,-14432.,-4468.7,-14620.,-16619.
142.0000000000,-18270.,-14337.,-4441.3,-14620.,-16619.
143.0000000000,-18147.,-14242.,-4414.3,-14620.,-16618.
144.0000000000,-18034.,-14157.,-4393.1,-14620.,-16618.
145.0000000000,-17917.,-14066.,-4367.2,-14620.,-16618.
146.0000000000,-17812.,-13986.,-4349.0,-14620.,-16617.
147.0000000000,-17698.,-13895.,-4322.7,-14619.,-16617.
148.0000000000,-17584.,-13805.,-4296.2,-14619.,-16616.
149.0000000000,-17471.,-13719.,-4271.5,-14619.,-16616.
150.0000000000,-17359.,-13632.,-4246.3,-14619.,-16616.
151.0000000000,-17248.,-13547.,-4221.7,-14619.,-16615.
152.0000000000,-17138.,-13463.,-4197.5,-14619.,-16615.
153.0000000000,-17030.,-13380.,-4173.9,-14619.,-16614.
154.0000000000,-16924.,-13299.,-4151.0,-14618.,-16614.
155.0000000000,-16818.,-13219.,-4128.2,-14618.,-16613.
156.0000000000,-16714.,-13140.,-4105.9,-14618.,-16613.
157.0000000000,-16612.,-13061.,-4083.9,-14618.,-16613.
158.0000000000,-16510.,-12985.,-4062.4,-14618.,-16612.
159.0000000000,-16413.,-12911.,-4042.9,-14618.,-16612.
160.0000000000,-16315.,-12836.,-4021.9,-14618.,-16611.
161.0000000000,-16218.,-12762.,-4001.1,-14618.,-16611.
162.0000000000,-16122.,-12688.,-3980.6,-14617.,-16611.
163.0000000000,-16026.,-12616.,-3960.4,-14617.,-16610.
164.0000000000,-15933.,-12545.,-3940.6,-14617.,-16610.
165.0000000000,-15841.,-12476.,-3922.2,-14617.,-16609.
166.0000000000,-15766.,-12422.,-3913.0,-14617.,-16609.
167.0000000000,-15680.,-12352.,-3894.1,-14617.,-16609.
168.0000000000,-15592.,-12282.,-3874.0,-14617.,-16608.
169.0000000000,-15504.,-12215.,-3854.9,-14616.,-16608.
170.0000000000,-15417.,-12148.,-3835.9,-14616.,-16607.
171.0000000000,-15331.,-12082.,-3817.1,-14616.,-16607.
172.0000000000,-15245.,-12017.,-3798.8,-14616.,-16606.
173.0000000000,-15161.,-11953.,-3780.8,-14616.,-16606.
174.0000000000,-15077.,-11890.,-3763.2,-14616.,-16606.
175.0000000000,-14995.,-11827.,-3745.9,-14616.,-16605.
176.0000000000,-14913.,-11766.,-3728.9,-14615.,-16605.
177.0000000000,-14833.,-11705.,-3712.1,-14615.,-16604.
178.0000000000,-14754.,-11645.,-3695.7,-14615.,-16604.
179.0000000000,-14675.,-11586.,-3679.4,-14615.,-16604.
180.0000000000,-14597.,-11527.,-3663.5,-14615.,-16603.
181.0000000000,-14524.,-11473.,-3650.1,-14615.,-16603.
182.0000000000,-14450.,-11416.,-3634.4,-14615.,-16602.
183.0000000000,-14376.,-11360.,-3619.3,-14614.,-16602.
184.0000000000,-14302.,-11303.,-3603.9,-14614.,-16602.
185.0000000000,-14229.,-11248.,-3588.7,-14614.,-16601.
186.0000000000,-14156.,-11193.,-3573.7,-14614.,-16601.
187.0000000000,-14085.,-11139.,-3559.0,-14614.,-16600.
188.0000000000,-14014.,-11086.,-3544.5,-14614.,-16600.
189.0000000000,-13944.,-11033.,-3530.3,-14614.,-16600.
190.0000000000,-13875.,-10981.,-3516.2,-14613.,-16599.
191.0000000000,-13806.,-10930.,-3502.3,-14613.,-16599.
192.0000000000,-13739.,-10879.,-3488.6,-14613.,-16598.
193.0000000000,-13672.,-10829.,-3475.1,-14613.,-16598.
194.0000000000,-13606.,-10779.,-3461.8,-14613.,-16598.
195.0000000000,-13541.,-10730.,-3448.6,-14613.,-16597.
196.0000000000,-13477.,-10683.,-3436.1,-14613.,-16597.
197.0000000000,-13422.,-10644.,-3429.3,-14613.,-16596.
198.0000000000,-13366.,-10600.,-3419.4,-14612.,-16596.
199.0000000000,-13306.,-10553.,-3406.4,-14612.,-16596.
200.0000000000,-13246.,-10506.,-3393.8,-14612.,-16595.
201.0000000000,-13185.,-10459.,-3380.5,-14612.,-16595.
202.0000000000,-13125.,-10413.,-3367.6,-14612.,-16594.
203.0000000000,-13065.,-10367.,-3355.2,-14612.,-16594.
204.0000000000,-13005.,-10322.,-3342.7,-14612.,-16594.
205.0000000000,-12946.,-10278.,-3330.5,-14612.,-16593.
206.0000000000,-12888.,-10234.,-3318.5,-14611.,-16593.
207.0000000000,-12830.,-10191.,-3306.8,-14611.,-16593.
208.0000000000,-12774.,-10149.,-3295.4,-14611.,-16592.
209.0000000000,-12717.,-10106.,-3284.0,-14611.,-16592.
210.0000000000,-12663.,-10066.,-3273.6,-14611.,-16591.
211.0000000000,-12608.,-10024.,-3262.5,-14611.,-16591.
212.0000000000,-12553.,-9983.3,-3251.4,-14611.,-16591.
213.0000000000,-12499.,-9942.8,-3240.5,-14611.,-16590.
214.0000000000,-12446.,-9902.8,-3229.8,-14610.,-16590.
215.0000000000,-12393.,-9863.3,-3219.2,-14610.,-16590.
216.0000000000,-12341.,-9824.2,-3208.7,-14610.,-16589.
217.0000000000,-12289.,-9785.5,-3198.4,-14610.,-16589.
218.0000000000,-12238.,-9747.2,-3188.2,-14610.,-16589.
219.0000000000,-12187.,-9709.4,-3178.1,-14610.,-16588.
220.0000000000,-12137.,-9671.9,-3168.2,-14610.,-16588.
221.0000000000,-12087.,-9634.9,-3158.3,-14610.,-16587.
222.0000000000,-12038.,-9598.2,-3148.6,-14609.,-16587.
223.0000000000,-11989.,-9562.0,-3139.0,-14609.,-16587.
224.0000000000,-11942.,-9526.5,-3129.8,-14609.,-16586.
225.0000000000,-11894.,-9490.9,-3120.4,-14609.,-16586.
226.0000000000,-11847.,-9455.6,-3111.0,-14609.,-16586.
227.0000000000,-11800.,-9420.7,-3101.8,-14609.,-16585.
228.0000000000,-11754.,-9386.2,-3092.7,-14609.,-16585.
229.0000000000,-11708.,-9352.1,-3083.6,-14609.,-16585.
230.0000000000,-11663.,-9318.3,-3074.7,-14609.,-16584.
231.0000000000,-11618.,-9284.9,-3065.9,-14608.,-16584.
232.0000000000,-11573.,-9251.7,-3057.2,-14608.,-16584.
233.0000000000,-11529.,-9219.0,-3048.5,-14608.,-16583.
234.0000000000,-11486.,-9186.8,-3040.1,-14608.,-16583.
235.0000000000,-11443.,-9154.6,-3031.7,-14608.,-16582.
236.0000000000,-11407.,-9129.7,-3027.8,-14608.,-16582.
237.0000000000,-11366.,-9097.6,-3019.4,-14608.,-16582.
238.0000000000,-11326.,-9066.4,-3011.2,-14608.,-16581.
239.0000000000,-11293.,-9043.7,-3008.3,-14608.,-16581.
240.0000000000,-11261.,-9018.8,-3004.3,-14607.,-16581.
241.0000000000,-11223.,-8986.0,-2994.9,-14607.,-16580.
242.0000000000,-11182.,-8953.7,-2985.5,-14607.,-16580.
243.0000000000,-11142.,-8922.4,-2976.3,-14607.,-16580.
244.0000000000,-11101.,-8891.8,-2967.5,-14607.,-16579.
245.0000000000,-11061.,-8861.8,-2959.1,-14607.,-16579.
246.0000000000,-11025.,-8835.4,-2952.8,-14607.,-16579.
247.0000000000,-10987.,-8806.0,-2944.7,-14607.,-16578.
248.0000000000,-10951.,-8779.2,-2938.1,-14607.,-16578.
249.0000000000,-10914.,-8751.7,-2931.0,-14606.,-16578.
250.0000000000,-10877.,-8722.9,-2923.0,-14606.,-16577.
251.0000000000,-10840.,-8694.5,-2915.0,-14606.,-16577.
252.0000000000,-10804.,-8668.6,-2908.6,-14606.,-16577.
253.0000000000,-10768.,-8641.2,-2901.1,-14606.,-16576.
254.0000000000,-10732.,-8614.7,-2894.2,-14606.,-16576.
255.0000000000,-10696.,-8587.5,-2886.7,-14606.,-16576.
256.0000000000,-10661.,-8560.7,-2879.3,-14606.,-16575.
257.0000000000,-10625.,-8534.2,-2872.0,-14606.,-16575.
258.0000000000,-10590.,-8508.0,-2864.9,-14606.,-16575.
259.0000000000,-10555.,-8482.2,-2857.9,-14605.,-16574.
260.0000000000,-10522.,-8458.2,-2852.0,-14605.,-16574.
261.0000000000,-10491.,-8436.0,-2847.3,-14605.,-16574.
262.0000000000,-10458.,-8411.2,-2840.8,-14605.,-16573.
263.0000000000,-10443.,-8405.0,-2846.4,-14605.,-16573.
264.0000000000,-10430.,-8393.7,-2849.2,-14605.,-16573.
265.0000000000,-10402.,-8364.7,-2840.3,-14605.,-16572.
266.0000000000,-10370.,-8336.2,-2830.9,-14605.,-16572.
267.0000000000,-10336.,-8309.2,-2822.0,-14605.,-16572.
268.0000000000,-10303.,-8283.3,-2813.8,-14605.,-16571.
269.0000000000,-10270.,-8258.2,-2806.0,-14604.,-16571.
270.0000000000,-10237.,-8233.7,-2798.6,-14604.,-16571.
271.0000000000,-10205.,-8209.6,-2791.5,-14604.,-16570.
272.0000000000,-10175.,-8188.6,-2786.3,-14604.,-16570.
273.0000000000,-10144.,-8165.1,-2779.5,-14604.,-16570.
274.0000000000,-10113.,-8141.7,-2772.7,-14604.,-16569.
275.0000000000,-10082.,-8118.7,-2766.2,-14604.,-16569.
276.0000000000,-10052.,-8096.1,-2759.8,-14604.,-16569.
277.0000000000,-10021.,-8073.8,-2753.5,-14604.,-16568.
278.0000000000,-9990.9,-8051.8,-2747.4,-14603.,-16568.
279.0000000000,-9961.1,-8030.0,-2741.3,-14603.,-16568.
280.0000000000,-9931.5,-8008.4,-2735.4,-14603.,-16567.
281.0000000000,-9902.2,-7987.0,-2729.6,-14603.,-16567.
282.0000000000,-9873.1,-7965.9,-2723.8,-14603.,-16567.
283.0000000000,-9844.3,-7944.9,-2718.1,-14603.,-16566.
284.0000000000,-9815.7,-7924.2,-2712.5,-14603.,-16566.
285.0000000000,-9787.4,-7903.6,-2706.9,-14603.,-16566.
286.0000000000,-9759.4,-7883.3,-2701.5,-14603.,-16565.
287.0000000000,-9733.8,-7865.4,-2697.5,-14603.,-16565.
288.0000000000,-9710.7,-7849.4,-2694.8,-14602.,-16565.
289.0000000000,-9696.5,-7841.5,-2697.5,-14602.,-16564.
290.0000000000,-9673.3,-7820.1,-2691.6,-14602.,-16564.
291.0000000000,-9647.0,-7798.2,-2684.9,-14602.,-16564.
292.0000000000,-9620.0,-7777.2,-2678.5,-14602.,-16563.
293.0000000000,-9593.0,-7756.8,-2672.3,-14602.,-16563.
294.0000000000,-9566.2,-7736.9,-2666.4,-14602.,-16563.
295.0000000000,-9539.6,-7717.4,-2660.7,-14602.,-16562.
296.0000000000,-9513.4,-7698.2,-2655.2,-14602.,-16562.
297.0000000000,-9487.4,-7679.2,-2649.8,-14602.,-16562.
298.0000000000,-9461.6,-7660.5,-2644.5,-14601.,-16561.
299.0000000000,-9436.1,-7642.0,-2639.4,-14601.,-16561.
300.0000000000,-9410.8,-7623.7,-2634.3,-14601.,-16561.
301.0000000000,-9385.8,-7605.6,-2629.3,-14601.,-16560.
302.0000000000,-9361.0,-7587.6,-2624.4,-14601.,-16560.
303.0000000000,-9336.4,-7569.9,-2619.5,-14601.,-16560.
304.0000000000,-9312.1,-7552.4,-2614.8,-14601.,-16559.
305.0000000000,-9287.9,-7534.9,-2610.0,-14601.,-16559.
306.0000000000,-9263.9,-7517.6,-2605.3,-14601.,-16559.
307.0000000000,-9240.2,-7500.4,-2600.7,-14601.,-16558.
308.0000000000,-9218.1,-7485.1,-2597.2,-14600.,-16558.
309.0000000000,-9195.5,-7468.5,-2592.9,-14600.,-16558.
310.0000000000,-9173.8,-7452.9,-2589.1,-14600.,-16557.
311.0000000000,-9152.2,-7437.1,-2585.2,-14600.,-16557.
312.0000000000,-9129.7,-7420.2,-2580.5,-14600.,-16557.
313.0000000000,-9108.2,-7404.8,-2576.7,-14600.,-16556.
314.0000000000,-9086.0,-7388.2,-2572.1,-14600.,-16556.
315.0000000000,-9063.7,-7371.7,-2567.5,-14600.,-16556.
316.0000000000,-9041.7,-7355.8,-2563.1,-14600.,-16555.
317.0000000000,-9019.8,-7339.8,-2558.7,-14600.,-16555.
318.0000000000,-8997.9,-7324.0,-2554.3,-14599.,-16555.
319.0000000000,-8976.2,-7308.3,-2550.0,-14599.,-16554.
320.0000000000,-8954.7,-7292.8,-2545.8,-14599.,-16554.
321.0000000000,-8933.3,-7277.4,-2541.6,-14599.,-16554.
322.0000000000,-8912.2,-7262.1,-2537.4,-14599.,-16553.
323.0000000000,-8891.2,-7247.0,-2533.3,-14599.,-16553.
324.0000000000,-8870.3,-7232.0,-2529.2,-14599.,-16553.
325.0000000000,-8849.7,-7217.2,-2525.2,-14599.,-16553.
326.0000000000,-8829.6,-7202.9,-2521.6,-14599.,-16552.
327.0000000000,-8809.9,-7188.8,-2517.9,-14598.,-16552.
328.0000000000,-8792.9,-7177.4,-2516.1,-14598.,-16552.
329.0000000000,-8776.1,-7165.2,-2513.8,-14598.,-16551.
330.0000000000,-8757.2,-7150.2,-2509.6,-14598.,-16551.
331.0000000000,-8737.5,-7135.3,-2505.3,-14598.,-16551.
332.0000000000,-8717.8,-7120.7,-2501.1,-14598.,-16550.
333.0000000000,-8698.1,-7106.3,-2497.0,-14598.,-16550.
334.0000000000,-8678.7,-7092.2,-2493.0,-14598.,-16550.
335.0000000000,-8659.3,-7078.3,-2489.1,-14598.,-16549.
336.0000000000,-8640.2,-7064.5,-2485.2,-14598.,-16549.
337.0000000000,-8621.2,-7050.8,-2481.4,-14597.,-16549.
338.0000000000,-8602.3,-7037.3,-2477.7,-14597.,-16548.
339.0000000000,-8583.6,-7023.8,-2474.0,-14597.,-16548.
340.0000000000,-8565.7,-7011.2,-2470.8,-14597.,-16548.
341.0000000000,-8547.4,-6997.9,-2467.1,-14597.,-16547.
342.0000000000,-8529.2,-6984.7,-2463.5,-14597.,-16547.
343.0000000000,-8511.0,-6971.7,-2459.9,-14597.,-16547.
344.0000000000,-8493.0,-6958.8,-2456.4,-14597.,-16546.
345.0000000000,-8475.1,-6946.0,-2452.9,-14597.,-16546.
346.0000000000,-8457.4,-6933.2,-2449.4,-14597.,-16546.
347.0000000000,-8439.8,-6920.6,-2446.0,-14596.,-16545.
348.0000000000,-8422.3,-6908.1,-2442.6,-14596.,-16545.
349.0000000000,-8404.9,-6895.7,-2439.2,-14596.,-16545.
350.0000000000,-8387.7,-6883.3,-2435.9,-14596.,-16544.
351.0000000000,-8370.6,-6871.1,-2432.6,-14596.,-16544.
352.0000000000,-8353.6,-6859.0,-2429.3,-14596.,-16544.
353.0000000000,-8336.7,-6846.9,-2426.0,-14596.,-16544.
354.0000000000,-8320.0,-6834.9,-2422.8,-14596.,-16543.
355.0000000000,-8305.6,-6825.4,-2421.1,-14596.,-16543.
356.0000000000,-8290.5,-6814.2,-2418.4,-14595.,-16543.
357.0000000000,-8274.5,-6802.1,-2415.1,-14595.,-16542.
358.0000000000,-8258.2,-6790.1,-2411.7,-14595.,-16542.
359.0000000000,-8242.0,-6778.2,-2408.3,-14595.,-16542.
360.0000000000,-8226.5,-6767.3,-2405.6,-14595.,-16542.
361.0000000000,-8212.2,-6757.3,-2403.4,-14595.,-16541.
362.0000000000,-8198.0,-6747.0,-2401.0,-14595.,-16541.
363.0000000000,-8182.6,-6735.2,-2397.7,-14595.,-16541.
364.0000000000,-8167.0,-6723.5,-2394.3,-14594.,-16541.
365.0000000000,-8151.3,-6712.1,-2391.0,-14594.,-16541.
366.0000000000,-8135.7,-6700.8,-2387.8,-14594.,-16541.
367.0000000000,-8120.3,-6689.7,-2384.7,-14594.,-16541.
368.0000000000,-8104.9,-6678.6,-2381.6,-14594.,-16540.
369.0000000000,-8089.7,-6667.7,-2378.6,-14594.,-16540.
370.0000000000,-8074.6,-6656.9,-2375.5,-14594.,-16540.
371.0000000000,-8059.6,-6646.1,-2372.6,-14593.,-16540.
372.0000000000,-8044.7,-6635.5,-2369.6,-14593.,-16540.
373.0000000000,-8029.9,-6624.9,-2366.7,-14593.,-16540.
374.0000000000,-8015.2,-6614.4,-2363.8,-14593.,-16540.
375.0000000000,-8000.6,-6604.0,-2361.0,-14593.,-16539.
376.0000000000,-7986.1,-6593.6,-2358.1,-14593.,-16539.
377.0000000000,-7971.7,-6583.3,-2355.3,-14593.,-16539.
378.0000000000,-7957.4,-6573.1,-2352.6,-14593.,-16539.
379.0000000000,-7943.2,-6563.0,-2349.8,-14592.,-16539.
380.0000000000,-7929.1,-6552.9,-2347.0,-14592.,-16539.
381.0000000000,-7915.1,-6542.9,-2344.3,-14592.,-16538.
382.0000000000,-7901.2,-6533.0,-2341.6,-14592.,-16538.
383.0000000000,-7887.4,-6523.1,-2338.9,-14592.,-16538.
384.0000000000,-7873.6,-6513.3,-2336.2,-14592.,-16538.
385.0000000000,-7860.0,-6503.6,-2333.6,-14592.,-16538.
386.0000000000,-7846.4,-6493.9,-2331.0,-14591.,-16537.
387.0000000000,-7833.0,-6484.3,-2328.3,-14591.,-16537.
388.0000000000,-7819.6,-6474.8,-2325.7,-14591.,-16537.
389.0000000000,-7806.5,-6465.5,-2323.3,-14591.,-16537.
390.0000000000,-7793.3,-6456.1,-2320.7,-14591.,-16537.
391.0000000000,-7780.2,-6446.7,-2318.2,-14591.,-16537.
392.0000000000,-7767.2,-6437.4,-2315.6,-14591.,-16536.
393.0000000000,-7754.3,-6428.1,-2313.1,-14590.,-16536.
394.0000000000,-7741.4,-6418.9,-2310.6,-14590.,-16536.
395.0000000000,-7728.6,-6409.8,-2308.1,-14590.,-16536.
396.0000000000,-7715.9,-6400.7,-2305.6,-14590.,-16536.
397.0000000000,-7703.3,-6391.7,-2303.1,-14590.,-16535.
398.0000000000,-7690.7,-6382.8,-2300.7,-14590.,-16535.
399.0000000000,-7678.3,-6373.9,-2298.3,-14590.,-16535.
400.0000000000,-7665.9,-6365.1,-2295.9,-14589.,-16535.
401.0000000000,-7653.6,-6356.3,-2293.5,-14589.,-16535.
402.0000000000,-7641.4,-6347.6,-2291.1,-14589.,-16534.
403.0000000000,-7629.2,-6338.9,-2288.7,-14589.,-16534.
404.0000000000,-7617.1,-6330.3,-2286.4,-14589.,-16534.
405.0000000000,-7605.1,-6321.8,-2284.0,-14589.,-16534.
406.0000000000,-7593.2,-6313.3,-2281.7,-14589.,-16534.
407.0000000000,-7581.3,-6304.8,-2279.4,-14588.,-16533.
408.0000000000,-7569.6,-6296.4,-2277.1,-14588.,-16533.
409.0000000000,-7557.9,-6288.1,-2274.8,-14588.,-16533.
410.0000000000,-7546.2,-6279.8,-2272.5,-14588.,-16533.
411.0000000000,-7534.6,-6271.6,-2270.3,-14588.,-16532.
412.0000000000,-7523.2,-6263.4,-2268.0,-14588.,-16532.
413.0000000000,-7511.7,-6255.2,-2265.8,-14588.,-16532.
414.0000000000,-7500.4,-6247.2,-2263.6,-14588.,-16532.
415.0000000000,-7489.1,-6239.1,-2261.3,-14587.,-16532.
416.0000000000,-7477.8,-6231.1,-2259.1,-14587.,-16531.
417.0000000000,-7466.7,-6223.2,-2257.0,-14587.,-16531.
418.0000000000,-7455.6,-6215.3,-2254.8,-14587.,-16531.
419.0000000000,-7444.6,-6207.5,-2252.6,-14587.,-16531.
420.0000000000,-7433.6,-6199.7,-2250.5,-14587.,-16530.
421.0000000000,-7422.8,-6192.1,-2248.4,-14587.,-16530.
422.0000000000,-7413.8,-6186.4,-2247.6,-14586.,-16530.
423.0000000000,-7404.2,-6179.1,-2245.9,-14586.,-16530.
424.0000000000,-7393.7,-6171.2,-2243.6,-14586.,-16530.
425.0000000000,-7383.1,-6163.3,-2241.3,-14586.,-16529.
426.0000000000,-7372.5,-6155.7,-2239.1,-14586.,-16529.
427.0000000000,-7361.9,-6148.0,-2236.9,-14586.,-16529.
428.0000000000,-7351.3,-6140.5,-2234.7,-14586.,-16529.
429.0000000000,-7340.9,-6133.0,-2232.6,-14585.,-16528.
430.0000000000,-7330.5,-6125.6,-2230.5,-14585.,-16528.
431.0000000000,-7320.1,-6118.3,-2228.4,-14585.,-16528.
432.0000000000,-7309.8,-6111.0,-2226.3,-14585.,-16528.
433.0000000000,-7299.6,-6103.7,-2224.3,-14585.,-16527.
434.0000000000,-7289.5,-6096.6,-2222.3,-14585.,-16527.
435.0000000000,-7279.5,-6089.4,-2220.3,-14585.,-16527.
436.0000000000,-7269.4,-6082.3,-2218.3,-14584.,-16527.
437.0000000000,-7259.4,-6075.3,-2216.3,-14584.,-16527.
438.0000000000,-7249.5,-6068.2,-2214.3,-14584.,-16526.
439.0000000000,-7239.6,-6061.3,-2212.4,-14584.,-16526.
440.0000000000,-7229.8,-6054.3,-2210.4,-14584.,-16526.
441.0000000000,-7220.1,-6047.4,-2208.5,-14584.,-16526.
442.0000000000,-7210.4,-6040.6,-2206.6,-14584.,-16525.
443.0000000000,-7200.7,-6033.8,-2204.7,-14583.,-16525.
444.0000000000,-7191.1,-6027.0,-2202.8,-14583.,-16525.
445.0000000000,-7181.6,-6020.3,-2200.9,-14583.,-16525.
446.0000000000,-7172.1,-6013.6,-2199.0,-14583.,-16524.
447.0000000000,-7162.6,-6006.9,-2197.1,-14583.,-16524.
448.0000000000,-7153.7,-6000.8,-2195.6,-14583.,-16524.
449.0000000000,-7144.4,-5994.1,-2193.7,-14583.,-16524.
450.0000000000,-7135.2,-5987.5,-2191.8,-14582.,-16523.
451.0000000000,-7126.0,-5981.1,-2190.0,-14582.,-16523.
452.0000000000,-7116.8,-5974.6,-2188.2,-14582.,-16523.
453.0000000000,-7107.7,-5968.1,-2186.3,-14582.,-16523.
454.0000000000,-7098.6,-5961.7,-2184.5,-14582.,-16522.
455.0000000000,-7089.5,-5955.3,-2182.7,-14582.,-16522.
456.0000000000,-7080.5,-5949.0,-2180.9,-14582.,-16522.
457.0000000000,-7071.6,-5942.7,-2179.1,-14581.,-16521.
458.0000000000,-7062.7,-5936.4,-2177.4,-14581.,-16521.
459.0000000000,-7055.3,-5931.9,-2176.7,-14581.,-16521.
460.0000000000,-7046.9,-5925.5,-2174.9,-14581.,-16521.
461.0000000000,-7038.3,-5919.2,-2173.1,-14581.,-16520.
462.0000000000,-7029.6,-5913.0,-2171.3,-14581.,-16520.
463.0000000000,-7021.1,-5906.9,-2169.5,-14581.,-16520.
464.0000000000,-7012.5,-5900.8,-2167.7,-14580.,-16520.
465.0000000000,-7003.8,-5894.7,-2166.0,-14580.,-16519.
466.0000000000,-6995.2,-5888.6,-2164.2,-14580.,-16519.
467.0000000000,-6986.7,-5882.6,-2162.5,-14580.,-16519.
468.0000000000,-6978.2,-5876.7,-2160.7,-14580.,-16519.
469.0000000000,-6969.8,-5870.8,-2159.0,-14580.,-16518.
470.0000000000,-6961.4,-5864.9,-2157.3,-14580.,-16518.
471.0000000000,-6953.1,-5859.0,-2155.7,-14579.,-16518.
472.0000000000,-6944.8,-5853.2,-2154.0,-14579.,-16518.
473.0000000000,-6936.5,-5847.5,-2152.3,-14579.,-16517.
474.0000000000,-6928.3,-5841.7,-2150.7,-14579.,-16517.
475.0000000000,-6920.3,-5836.2,-2149.2,-14579.,-16517.
476.0000000000,-6912.2,-5830.6,-2147.6,-14579.,-16516.
477.0000000000,-6904.1,-5824.9,-2145.9,-14579.,-16516.
478.0000000000,-6896.1,-5819.3,-2144.3,-14578.,-16516.
479.0000000000,-6888.0,-5813.7,-2142.7,-14578.,-16516.
480.0000000000,-6880.1,-5808.1,-2141.1,-14578.,-16515.
481.0000000000,-6872.1,-5802.6,-2139.5,-14578.,-16515.
482.0000000000,-6864.2,-5797.1,-2137.9,-14578.,-16515.
483.0000000000,-6856.4,-5791.7,-2136.4,-14578.,-16515.
484.0000000000,-6848.6,-5786.3,-2134.8,-14578.,-16514.
485.0000000000,-6840.8,-5780.9,-2133.2,-14577.,-16514.
486.0000000000,-6833.1,-5775.5,-2131.7,-14577.,-16514.
487.0000000000,-6825.4,-5770.2,-2130.2,-14577.,-16513.
488.0000000000,-6817.7,-5764.9,-2128.6,-14577.,-16513.
489.0000000000,-6810.1,-5759.6,-2127.1,-14577.,-16513.
490.0000000000,-6802.5,-5754.3,-2125.6,-14577.,-16513.
491.0000000000,-6795.0,-5749.1,-2124.1,-14576.,-16512.
492.0000000000,-6788.6,-5745.2,-2123.4,-14576.,-16512.
493.0000000000,-6781.5,-5739.9,-2121.9,-14576.,-16512.
494.0000000000,-6774.6,-5735.2,-2120.7,-14576.,-16511.
495.0000000000,-6768.4,-5731.0,-2119.8,-14576.,-16511.
496.0000000000,-6761.3,-5725.6,-2118.2,-14576.,-16511.
497.0000000000,-6754.1,-5720.3,-2116.6,-14576.,-16511.
498.0000000000,-6747.8,-5716.3,-2115.8,-14575.,-16510.
499.0000000000,-6741.0,-5711.3,-2114.4,-14575.,-16510.
500.0000000000,-6733.9,-5706.0,-2112.7,-14575.,-16510.
501.0000000000,-6726.7,-5700.8,-2111.1,-14575.,-16509.
502.0000000000,-6719.4,-5695.7,-2109.5,-14575.,-16509.
503.0000000000,-6712.2,-5690.7,-2107.9,-14575.,-16509.
504.0000000000,-6705.0,-5685.7,-2106.4,-14575.,-16509.
505.0000000000,-6697.9,-5680.8,-2104.9,-14574.,-16508.
506.0000000000,-6690.8,-5675.9,-2103.4,-14574.,-16508.
507.0000000000,-6683.8,-5671.0,-2101.9,-14574.,-16508.
508.0000000000,-6677.2,-5666.7,-2100.8,-14574.,-16507.
509.0000000000,-6670.4,-5661.8,-2099.4,-14574.,-16507.
510.0000000000,-6664.6,-5658.2,-2098.7,-14574.,-16507.
511.0000000000,-6665.0,-5661.2,-2102.4,-14573.,-16507.
512.0000000000,-6660.7,-5656.0,-2101.1,-14573.,-16506.
513.0000000000,-6654.5,-5650.0,-2098.9,-14573.,-16506.
514.0000000000,-6647.6,-5644.4,-2096.8,-14573.,-16506.
515.0000000000,-6640.5,-5639.1,-2094.9,-14573.,-16505.
516.0000000000,-6633.5,-5634.0,-2093.1,-14573.,-16505.
517.0000000000,-6626.5,-5629.0,-2091.4,-14573.,-16505.
518.0000000000,-6619.6,-5624.2,-2089.7,-14572.,-16504.
519.0000000000,-6612.8,-5619.4,-2088.1,-14572.,-16504.
520.0000000000,-6606.0,-5614.7,-2086.6,-14572.,-16504.
521.0000000000,-6599.2,-5610.0,-2085.1,-14572.,-16504.
522.0000000000,-6592.5,-5605.5,-2083.6,-14572.,-16503.
523.0000000000,-6585.9,-5600.9,-2082.1,-14572.,-16503.
524.0000000000,-6579.2,-5596.4,-2080.7,-14571.,-16503.
525.0000000000,-6572.8,-5592.0,-2079.4,-14571.,-16502.
526.0000000000,-6566.3,-5587.7,-2078.0,-14571.,-16502.
527.0000000000,-6559.8,-5583.2,-2076.7,-14571.,-16502.
528.0000000000,-6553.6,-5579.1,-2075.5,-14571.,-16502.
529.0000000000,-6548.6,-5576.3,-2075.1,-14571.,-16501.
530.0000000000,-6545.3,-5574.7,-2075.7,-14571.,-16501.
531.0000000000,-6539.8,-5569.9,-2074.2,-14570.,-16501.
532.0000000000,-6533.6,-5565.0,-2072.5,-14570.,-16500.
533.0000000000,-6527.2,-5560.4,-2070.9,-14570.,-16500.
534.0000000000,-6520.8,-5555.8,-2069.3,-14570.,-16500.
535.0000000000,-6514.4,-5551.4,-2067.8,-14570.,-16499.
536.0000000000,-6523.4,-5564.2,-2077.7,-14570.,-16499.
537.0000000000,-6528.1,-5565.6,-2080.8,-14569.,-16499.
538.0000000000,-6526.8,-5560.6,-2079.5,-14569.,-16499.
539.0000000000,-6521.5,-5553.3,-2076.3,-14569.,-16498.
540.0000000000,-6515.0,-5547.0,-2073.3,-14569.,-16498.
541.0000000000,-6513.7,-5547.4,-2074.7,-14569.,-16498.
542.0000000000,-6508.5,-5541.4,-2072.2,-14569.,-16497.
543.0000000000,-6502.0,-5535.4,-2069.5,-14569.,-16497.
544.0000000000,-6495.3,-5530.1,-2067.0,-14568.,-16497.
545.0000000000,-6488.5,-5524.9,-2064.8,-14568.,-16496.
546.0000000000,-6481.8,-5520.1,-2062.7,-14568.,-16496.
547.0000000000,-6475.2,-5515.4,-2060.7,-14568.,-16496.
548.0000000000,-6468.6,-5510.9,-2058.9,-14568.,-16496.
549.0000000000,-6462.2,-5506.5,-2057.2,-14568.,-16495.
550.0000000000,-6455.7,-5502.1,-2055.6,-14567.,-16495.
551.0000000000,-6449.4,-5497.9,-2054.0,-14567.,-16495.
552.0000000000,-6443.1,-5493.7,-2052.4,-14567.,-16494.
553.0000000000,-6436.9,-5489.6,-2051.0,-14567.,-16494.
554.0000000000,-6430.7,-5485.5,-2049.5,-14567.,-16494.
555.0000000000,-6424.5,-5481.5,-2048.1,-14567.,-16493.
556.0000000000,-6418.5,-5477.6,-2046.8,-14566.,-16493.
557.0000000000,-6412.5,-5473.7,-2045.5,-14566.,-16493.
558.0000000000,-6407.6,-5471.1,-2045.0,-14566.,-16492.
559.0000000000,-6402.0,-5467.1,-2043.7,-14566.,-16492.
560.0000000000,-6396.1,-5463.0,-2042.3,-14566.,-16492.
561.0000000000,-6390.1,-5459.0,-2040.9,-14566.,-16492.
562.0000000000,-6385.7,-5456.8,-2040.7,-14566.,-16491.
563.0000000000,-6382.1,-5454.9,-2040.7,-14565.,-16491.
564.0000000000,-6378.2,-5452.1,-2040.2,-14565.,-16491.
565.0000000000,-6372.8,-5447.8,-2038.7,-14565.,-16490.
566.0000000000,-6367.1,-5443.5,-2037.1,-14565.,-16490.
567.0000000000,-6361.2,-5439.4,-2035.5,-14565.,-16490.
568.0000000000,-6355.3,-5435.4,-2034.1,-14565.,-16489.
569.0000000000,-6349.4,-5431.5,-2032.7,-14564.,-16489.
570.0000000000,-6343.6,-5427.7,-2031.3,-14564.,-16489.
571.0000000000,-6338.5,-5424.7,-2030.5,-14564.,-16489.
572.0000000000,-6333.0,-5420.9,-2029.2,-14564.,-16488.
573.0000000000,-6327.3,-5417.1,-2027.9,-14564.,-16488.
574.0000000000,-6321.7,-5413.4,-2026.6,-14564.,-16488.
575.0000000000,-6316.1,-5409.8,-2025.4,-14563.,-16487.
576.0000000000,-6310.5,-5406.2,-2024.2,-14563.,-16487.
577.0000000000,-6304.9,-5402.6,-2023.0,-14563.,-16487.
578.0000000000,-6299.4,-5399.0,-2021.8,-14563.,-16486.
579.0000000000,-6296.5,-5398.5,-2022.6,-14563.,-16486.
580.0000000000,-6298.9,-5402.7,-2026.6,-14563.,-16486.
581.0000000000,-6295.7,-5398.0,-2025.1,-14563.,-16485.
582.0000000000,-6290.7,-5393.1,-2023.1,-14562.,-16485.
583.0000000000,-6285.1,-5388.7,-2021.3,-14562.,-16485.
584.0000000000,-6279.5,-5384.5,-2019.6,-14562.,-16484.
585.0000000000,-6273.8,-5380.6,-2018.0,-14562.,-16484.
586.0000000000,-6268.2,-5376.8,-2016.5,-14562.,-16484.
587.0000000000,-6262.7,-5373.1,-2015.1,-14562.,-16484.
588.0000000000,-6257.2,-5369.5,-2013.8,-14561.,-16483.
589.0000000000,-6252.4,-5366.8,-2013.0,-14561.,-16483.
590.0000000000,-6248.9,-5365.1,-2013.0,-14561.,-16483.
591.0000000000,-6244.1,-5361.4,-2011.7,-14561.,-16482.
592.0000000000,-6238.9,-5357.6,-2010.3,-14561.,-16482.
593.0000000000,-6233.6,-5354.0,-2008.9,-14561.,-16482.
594.0000000000,-6228.6,-5351.0,-2008.0,-14560.,-16481.
595.0000000000,-6225.6,-5349.9,-2008.3,-14560.,-16481.
596.0000000000,-6223.6,-5349.2,-2009.0,-14560.,-16481.
597.0000000000,-6219.3,-5345.2,-2007.5,-14560.,-16480.
598.0000000000,-6214.2,-5341.2,-2005.9,-14560.,-16480.
599.0000000000,-6209.0,-5337.4,-2004.4,-14560.,-16480.
600.0000000000,-6203.7,-5333.8,-2003.0,-14559.,-16480.
601.0000000000,-6198.4,-5330.3,-2001.7,-14559.,-16479.
602.0000000000,-6193.2,-5326.9,-2000.4,-14559.,-16479.
603.0000000000,-6188.0,-5323.5,-1999.2,-14559.,-16479.
604.0000000000,-6182.8,-5320.2,-1998.0,-14559.,-16478.
605.0000000000,-6177.8,-5317.1,-1996.9,-14559.,-16478.
606.0000000000,-6172.7,-5313.8,-1995.7,-14558.,-16478.
607.0000000000,-6168.0,-5311.0,-1994.9,-14558.,-16477.
608.0000000000,-6163.2,-5307.9,-1993.8,-14558.,-16477.
609.0000000000,-6158.2,-5304.7,-1992.7,-14558.,-16477.
610.0000000000,-6153.3,-5301.6,-1991.6,-14558.,-16476.
611.0000000000,-6148.3,-5298.5,-1990.6,-14558.,-16476.
612.0000000000,-6143.4,-5295.4,-1989.5,-14557.,-16476.
613.0000000000,-6140.7,-5294.8,-1990.1,-14557.,-16475.
614.0000000000,-6137.0,-5292.2,-1989.4,-14557.,-16475.
615.0000000000,-6132.5,-5288.8,-1988.2,-14557.,-16475.
616.0000000000,-6129.3,-5287.2,-1988.2,-14557.,-16474.
617.0000000000,-6124.9,-5283.8,-1987.0,-14557.,-16474.
618.0000000000,-6120.1,-5280.4,-1985.7,-14556.,-16474.
619.0000000000,-6115.3,-5277.1,-1984.4,-14556.,-16474.
620.0000000000,-6110.5,-5274.0,-1983.3,-14556.,-16473.
621.0000000000,-6106.3,-5271.6,-1982.6,-14556.,-16473.
622.0000000000,-6102.2,-5269.1,-1981.9,-14556.,-16473.
623.0000000000,-6097.6,-5266.0,-1980.8,-14556.,-16472.
624.0000000000,-6093.0,-5262.8,-1979.6,-14555.,-16472.
625.0000000000,-6088.6,-5260.2,-1978.8,-14555.,-16472.
626.0000000000,-6084.0,-5257.2,-1977.7,-14555.,-16471.
627.0000000000,-6083.0,-5258.3,-1979.4,-14555.,-16471.
628.0000000000,-6079.8,-5255.3,-1978.5,-14555.,-16471.
629.0000000000,-6077.3,-5253.8,-1978.5,-14555.,-16470.
630.0000000000,-6074.2,-5251.5,-1977.9,-14554.,-16470.
631.0000000000,-6069.9,-5247.9,-1976.5,-14554.,-16470.
632.0000000000,-6065.3,-5244.4,-1975.1,-14554.,-16469.
633.0000000000,-6060.6,-5241.2,-1973.7,-14554.,-16469.
634.0000000000,-6056.0,-5238.2,-1972.5,-14554.,-16469.
635.0000000000,-6059.3,-5244.2,-1977.3,-14554.,-16468.
636.0000000000,-6058.5,-5242.0,-1977.1,-14553.,-16468.
637.0000000000,-6054.8,-5237.6,-1975.2,-14553.,-16468.
638.0000000000,-6050.2,-5233.6,-1973.4,-14553.,-16468.
639.0000000000,-6045.4,-5229.9,-1971.7,-14553.,-16467.
640.0000000000,-6040.6,-5226.5,-1970.2,-14553.,-16467.
641.0000000000,-6035.8,-5223.2,-1968.8,-14553.,-16467.
642.0000000000,-6031.0,-5220.1,-1967.4,-14552.,-16466.
643.0000000000,-6026.3,-5217.1,-1966.2,-14552.,-16466.
644.0000000000,-6021.7,-5214.2,-1965.0,-14552.,-16466.
645.0000000000,-6017.1,-5211.3,-1963.9,-14552.,-16465.
646.0000000000,-6012.6,-5208.5,-1962.8,-14552.,-16465.
647.0000000000,-6008.0,-5205.7,-1961.7,-14552.,-16465.
648.0000000000,-6003.6,-5202.9,-1960.7,-14551.,-16464.
649.0000000000,-6002.4,-5203.9,-1962.1,-14551.,-16464.
650.0000000000,-5999.0,-5200.9,-1961.1,-14551.,-16464.
651.0000000000,-5994.8,-5197.7,-1959.8,-14551.,-16463.
652.0000000000,-5990.4,-5194.6,-1958.6,-14551.,-16463.
653.0000000000,-5985.9,-5191.7,-1957.4,-14551.,-16463.
654.0000000000,-5981.5,-5188.9,-1956.3,-14550.,-16462.
655.0000000000,-5977.1,-5186.2,-1955.3,-14550.,-16462.
656.0000000000,-5972.7,-5183.4,-1954.2,-14550.,-16462.
657.0000000000,-5968.3,-5180.8,-1953.2,-14550.,-16462.
658.0000000000,-5964.0,-5178.2,-1952.3,-14550.,-16461.
659.0000000000,-5959.9,-5175.7,-1951.4,-14550.,-16461.
660.0000000000,-5956.3,-5173.8,-1951.0,-14549.,-16461.
661.0000000000,-5954.1,-5173.3,-1951.4,-14549.,-16460.
662.0000000000,-5950.5,-5170.5,-1950.4,-14549.,-16460.
663.0000000000,-5946.4,-5167.5,-1949.3,-14549.,-16460.
664.0000000000,-5942.2,-5164.8,-1948.2,-14549.,-16459.
665.0000000000,-5938.0,-5162.1,-1947.2,-14549.,-16459.
666.0000000000,-5933.8,-5159.4,-1946.2,-14548.,-16459.
667.0000000000,-5929.6,-5156.9,-1945.2,-14548.,-16458.
668.0000000000,-5925.4,-5154.3,-1944.3,-14548.,-16458.
669.0000000000,-5921.3,-5151.8,-1943.4,-14548.,-16458.
670.0000000000,-5917.2,-5149.3,-1942.5,-14548.,-16457.
671.0000000000,-5913.1,-5146.9,-1941.6,-14547.,-16457.
672.0000000000,-5909.0,-5144.4,-1940.7,-14547.,-16457.
673.0000000000,-5905.0,-5142.0,-1939.9,-14547.,-16456.
674.0000000000,-5912.0,-5152.2,-1947.3,-14547.,-16456.
675.0000000000,-5917.4,-5155.6,-1950.9,-14547.,-16456.
676.0000000000,-5916.2,-5151.0,-1949.1,-14547.,-16455.
677.0000000000,-5912.7,-5146.5,-1946.9,-14546.,-16455.
678.0000000000,-5908.4,-5142.5,-1944.9,-14546.,-16455.
679.0000000000,-5903.9,-5138.9,-1943.0,-14546.,-16454.
680.0000000000,-5899.5,-5135.6,-1941.4,-14546.,-16454.
681.0000000000,-5895.1,-5132.6,-1939.9,-14546.,-16454.
682.0000000000,-5890.7,-5129.7,-1938.6,-14546.,-16453.
683.0000000000,-5886.4,-5127.0,-1937.3,-14545.,-16453.
684.0000000000,-5882.2,-5124.3,-1936.1,-14545.,-16453.
685.0000000000,-5878.0,-5121.7,-1935.0,-14545.,-16453.
686.0000000000,-5873.9,-5119.1,-1933.9,-14545.,-16452.
687.0000000000,-5869.8,-5116.6,-1932.9,-14545.,-16452.
688.0000000000,-5865.8,-5114.2,-1931.9,-14545.,-16452.
689.0000000000,-5861.7,-5111.8,-1930.9,-14544.,-16451.
690.0000000000,-5857.7,-5109.4,-1930.0,-14544.,-16451.
691.0000000000,-5853.8,-5107.0,-1929.1,-14544.,-16451.
692.0000000000,-5850.8,-5105.8,-1929.0,-14544.,-16450.
693.0000000000,-5847.2,-5103.4,-1928.1,-14544.,-16450.
694.0000000000,-5843.4,-5100.9,-1927.1,-14543.,-16450.
695.0000000000,-5839.5,-5098.5,-1926.2,-14543.,-16449.
696.0000000000,-5835.6,-5096.2,-1925.3,-14543.,-16449.
697.0000000000,-5831.7,-5093.9,-1924.4,-14543.,-16449.
698.0000000000,-5827.9,-5091.6,-1923.5,-14543.,-16448.
699.0000000000,-5824.0,-5089.3,-1922.7,-14543.,-16448.
700.0000000000,-5820.2,-5087.1,-1921.9,-14542.,-16448.
701.0000000000,-5816.5,-5084.9,-1921.1,-14542.,-16447.
702.0000000000,-5812.7,-5082.6,-1920.3,-14542.,-16447.
703.0000000000,-5809.0,-5080.5,-1919.5,-14542.,-16447.
704.0000000000,-5805.2,-5078.3,-1918.7,-14542.,-16446.
705.0000000000,-5801.5,-5076.1,-1917.9,-14542.,-16446.
706.0000000000,-5797.9,-5074.0,-1917.1,-14541.,-16446.
707.0000000000,-5794.2,-5071.8,-1916.4,-14541.,-16445.
708.0000000000,-5790.5,-5069.7,-1915.6,-14541.,-16445.
709.0000000000,-5786.9,-5067.6,-1914.9,-14541.,-16445.
710.0000000000,-5783.4,-5065.5,-1914.2,-14541.,-16444.
711.0000000000,-5779.8,-5063.4,-1913.4,-14540.,-16444.
712.0000000000,-5776.2,-5061.3,-1912.7,-14540.,-16444.
713.0000000000,-5772.6,-5059.2,-1911.9,-14540.,-16443.
714.0000000000,-5769.1,-5057.1,-1911.2,-14540.,-16443.
715.0000000000,-5765.5,-5055.1,-1910.5,-14540.,-16443.
716.0000000000,-5762.0,-5053.0,-1909.8,-14540.,-16443.
717.0000000000,-5758.5,-5050.9,-1909.0,-14539.,-16442.
718.0000000000,-5755.1,-5049.0,-1908.4,-14539.,-16442.
719.0000000000,-5751.7,-5047.0,-1907.7,-14539.,-16442.
720.0000000000,-5748.2,-5044.9,-1907.0,-14539.,-16441.
721.0000000000,-5744.8,-5042.9,-1906.3,-14539.,-16441.
722.0000000000,-5741.4,-5041.0,-1905.6,-14539.,-16441.
723.0000000000,-5738.2,-5039.1,-1905.0,-14538.,-16440.
724.0000000000,-5734.8,-5037.1,-1904.3,-14538.,-16440.
725.0000000000,-5731.4,-5035.1,-1903.6,-14538.,-16440.
726.0000000000,-5728.0,-5033.1,-1902.9,-14538.,-16439.
727.0000000000,-5728.8,-5035.9,-1905.4,-14538.,-16439.
728.0000000000,-5726.9,-5033.7,-1904.8,-14537.,-16439.
729.0000000000,-5723.9,-5031.0,-1903.7,-14537.,-16438.
730.0000000000,-5720.8,-5028.8,-1902.8,-14537.,-16438.
731.0000000000,-5718.2,-5027.4,-1902.4,-14537.,-16438.
732.0000000000,-5716.3,-5026.5,-1902.5,-14537.,-16437.
733.0000000000,-5714.7,-5025.7,-1902.6,-14537.,-16437.
734.0000000000,-5711.8,-5023.1,-1901.5,-14536.,-16437.
735.0000000000,-5708.4,-5020.6,-1900.4,-14536.,-16436.
736.0000000000,-5705.0,-5018.3,-1899.4,-14536.,-16436.
737.0000000000,-5701.5,-5016.0,-1898.4,-14536.,-16436.
738.0000000000,-5698.1,-5013.9,-1897.5,-14536.,-16435.
739.0000000000,-5694.8,-5011.9,-1896.7,-14535.,-16435.
740.0000000000,-5693.4,-5012.1,-1897.4,-14535.,-16435.
741.0000000000,-5690.9,-5010.1,-1896.7,-14535.,-16434.
742.0000000000,-5687.8,-5007.8,-1895.7,-14535.,-16434.
743.0000000000,-5684.4,-5005.5,-1894.8,-14535.,-16434.
744.0000000000,-5681.1,-5003.4,-1893.9,-14535.,-16433.
745.0000000000,-5677.7,-5001.3,-1893.0,-14534.,-16433.
746.0000000000,-5674.4,-4999.3,-1892.2,-14534.,-16433.
747.0000000000,-5671.1,-4997.3,-1891.4,-14534.,-16432.
748.0000000000,-5667.8,-4995.3,-1890.7,-14534.,-16432.
749.0000000000,-5664.5,-4993.4,-1889.9,-14534.,-16432.
750.0000000000,-5661.3,-4991.5,-1889.2,-14533.,-16431.
751.0000000000,-5658.0,-4989.6,-1888.5,-14533.,-16431.
752.0000000000,-5656.2,-4989.2,-1888.8,-14533.,-16431.
753.0000000000,-5654.9,-4989.0,-1889.2,-14533.,-16430.
754.0000000000,-5652.4,-4986.9,-1888.5,-14533.,-16430.
755.0000000000,-5649.3,-4984.6,-1887.5,-14533.,-16430.
756.0000000000,-5646.1,-4982.5,-1886.6,-14532.,-16430.
757.0000000000,-5642.9,-4980.4,-1885.8,-14532.,-16429.
758.0000000000,-5639.6,-4978.4,-1885.0,-14532.,-16429.
759.0000000000,-5636.4,-4976.5,-1884.2,-14532.,-16429.
760.0000000000,-5633.3,-4974.6,-1883.4,-14532.,-16428.
761.0000000000,-5631.3,-4974.1,-1883.6,-14531.,-16428.
762.0000000000,-5630.2,-4974.1,-1884.2,-14531.,-16428.
763.0000000000,-5627.7,-4971.9,-1883.3,-14531.,-16427.
764.0000000000,-5624.7,-4969.6,-1882.4,-14531.,-16427.
765.0000000000,-5621.6,-4967.6,-1881.6,-14531.,-16427.
766.0000000000,-5618.4,-4965.6,-1880.7,-14531.,-16426.
767.0000000000,-5615.3,-4963.6,-1879.9,-14530.,-16426.
768.0000000000,-5612.1,-4961.7,-1879.1,-14530.,-16426.
769.0000000000,-5609.0,-4959.8,-1878.4,-14530.,-16425.
770.0000000000,-5605.9,-4958.0,-1877.7,-14530.,-16425.
771.0000000000,-5602.8,-4956.1,-1877.0,-14530.,-16425.
772.0000000000,-5599.8,-4954.3,-1876.3,-14529.,-16424.
773.0000000000,-5596.7,-4952.5,-1875.6,-14529.,-16424.
774.0000000000,-5593.7,-4950.7,-1874.9,-14529.,-16424.
775.0000000000,-5590.7,-4948.9,-1874.3,-14529.,-16423.
776.0000000000,-5587.7,-4947.2,-1873.6,-14529.,-16423.
777.0000000000,-5584.7,-4945.5,-1873.0,-14529.,-16423.
778.0000000000,-5581.9,-4943.9,-1872.4,-14528.,-16422.
779.0000000000,-5578.9,-4942.1,-1871.8,-14528.,-16422.
780.0000000000,-5576.0,-4940.4,-1871.2,-14528.,-16422.
781.0000000000,-5573.1,-4938.6,-1870.5,-14528.,-16421.
782.0000000000,-5570.1,-4936.9,-1869.9,-14528.,-16421.
783.0000000000,-5567.2,-4935.2,-1869.3,-14527.,-16421.
784.0000000000,-5564.3,-4933.5,-1868.7,-14527.,-16420.
785.0000000000,-5561.4,-4931.8,-1868.1,-14527.,-16420.
786.0000000000,-5558.5,-4930.1,-1867.5,-14527.,-16420.
787.0000000000,-5555.6,-4928.4,-1866.9,-14527.,-16419.
788.0000000000,-5552.7,-4926.7,-1866.3,-14526.,-16419.
789.0000000000,-5550.4,-4925.6,-1866.0,-14526.,-16419.
790.0000000000,-5547.8,-4924.0,-1865.6,-14526.,-16418.
791.0000000000,-5545.1,-4922.3,-1865.0,-14526.,-16418.
792.0000000000,-5542.3,-4920.6,-1864.3,-14526.,-16418.
793.0000000000,-5539.5,-4918.9,-1863.7,-14526.,-16417.
794.0000000000,-5538.5,-4919.3,-1864.5,-14525.,-16417.
795.0000000000,-5536.2,-4917.4,-1863.8,-14525.,-16417.
796.0000000000,-5533.5,-4915.4,-1863.0,-14525.,-16416.
797.0000000000,-5531.3,-4914.2,-1862.8,-14525.,-16416.
798.0000000000,-5528.8,-4912.5,-1862.1,-14525.,-16416.
799.0000000000,-5526.2,-4911.0,-1861.6,-14524.,-16416.
800.0000000000,-5523.5,-4909.1,-1860.8,-14524.,-16415.
801.0000000000,-5520.7,-4907.3,-1860.1,-14524.,-16415.
802.0000000000,-5517.9,-4905.6,-1859.4,-14524.,-16415.
803.0000000000,-5515.0,-4903.8,-1858.8,-14524.,-16414.
804.0000000000,-5512.2,-4902.2,-1858.1,-14524.,-16414.
805.0000000000,-5509.5,-4900.5,-1857.5,-14523.,-16414.
806.0000000000,-5506.7,-4898.8,-1856.9,-14523.,-16413.
807.0000000000,-5504.3,-4897.7,-1856.6,-14523.,-16413.
808.0000000000,-5501.7,-4896.0,-1856.0,-14523.,-16413.
809.0000000000,-5501.1,-4896.7,-1856.9,-14523.,-16412.
810.0000000000,-5506.4,-4903.5,-1861.9,-14522.,-16412.
811.0000000000,-5510.3,-4905.6,-1864.3,-14522.,-16412.
812.0000000000,-5509.4,-4902.1,-1862.7,-14522.,-16411.
813.0000000000,-5506.8,-4898.8,-1861.0,-14522.,-16411.
814.0000000000,-5503.8,-4895.9,-1859.5,-14522.,-16411.
815.0000000000,-5500.9,-4893.7,-1858.3,-14521.,-16410.
816.0000000000,-5497.9,-4891.4,-1857.1,-14521.,-16410.
817.0000000000,-5494.8,-4889.2,-1856.0,-14521.,-16410.
818.0000000000,-5491.8,-4887.2,-1855.0,-14521.,-16409.
819.0000000000,-5488.9,-4885.3,-1854.0,-14521.,-16409.
820.0000000000,-5485.9,-4883.4,-1853.1,-14521.,-16409.
821.0000000000,-5483.0,-4881.6,-1852.3,-14520.,-16408.
822.0000000000,-5480.1,-4879.9,-1851.5,-14520.,-16408.
823.0000000000,-5477.3,-4878.2,-1850.8,-14520.,-16408.
824.0000000000,-5474.4,-4876.5,-1850.1,-14520.,-16407.
825.0000000000,-5471.6,-4874.8,-1849.4,-14520.,-16407.
826.0000000000,-5469.2,-4873.6,-1849.0,-14519.,-16407.
827.0000000000,-5466.5,-4871.9,-1848.3,-14519.,-16406.
828.0000000000,-5463.9,-4870.4,-1847.7,-14519.,-16406.
829.0000000000,-5462.1,-4869.8,-1847.7,-14519.,-16406.
830.0000000000,-5459.6,-4868.0,-1847.0,-14519.,-16405.
831.0000000000,-5456.9,-4866.3,-1846.3,-14518.,-16405.
832.0000000000,-5454.8,-4865.3,-1846.0,-14518.,-16405.
833.0000000000,-5455.5,-4867.4,-1847.8,-14518.,-16404.
834.0000000000,-5453.8,-4865.3,-1847.1,-14518.,-16404.
835.0000000000,-5451.3,-4863.2,-1846.1,-14518.,-16404.
836.0000000000,-5450.3,-4863.1,-1846.5,-14518.,-16403.
837.0000000000,-5448.4,-4861.6,-1845.9,-14517.,-16403.
838.0000000000,-5448.4,-4862.4,-1846.9,-14517.,-16403.
839.0000000000,-5446.4,-4860.3,-1845.9,-14517.,-16402.
840.0000000000,-5443.8,-4858.0,-1844.8,-14517.,-16402.
841.0000000000,-5441.0,-4855.9,-1843.8,-14517.,-16402.
842.0000000000,-5438.1,-4854.0,-1842.9,-14516.,-16402.
843.0000000000,-5435.3,-4852.2,-1842.0,-14516.,-16401.
844.0000000000,-5434.4,-4852.6,-1842.6,-14516.,-16401.
845.0000000000,-5432.1,-4850.7,-1841.8,-14516.,-16401.
846.0000000000,-5429.5,-4848.8,-1840.9,-14516.,-16400.
847.0000000000,-5429.8,-4850.6,-1842.5,-14515.,-16400.
848.0000000000,-5428.0,-4848.5,-1841.6,-14515.,-16400.
849.0000000000,-5425.5,-4846.3,-1840.6,-14515.,-16399.
850.0000000000,-5422.7,-4844.3,-1839.6,-14515.,-16399.
851.0000000000,-5419.9,-4842.5,-1838.7,-14515.,-16399.
852.0000000000,-5417.1,-4840.7,-1837.9,-14515.,-16398.
853.0000000000,-5414.4,-4839.1,-1837.1,-14514.,-16398.
854.0000000000,-5411.6,-4837.4,-1836.4,-14514.,-16398.
855.0000000000,-5409.0,-4835.9,-1835.7,-14514.,-16397.
856.0000000000,-5406.3,-4834.3,-1835.0,-14514.,-16397.
857.0000000000,-5403.7,-4832.9,-1834.4,-14514.,-16397.
858.0000000000,-5401.1,-4831.3,-1833.8,-14513.,-16396.
859.0000000000,-5398.4,-4829.8,-1833.1,-14513.,-16396.
860.0000000000,-5395.8,-4828.3,-1832.5,-14513.,-16396.
861.0000000000,-5402.8,-4838.0,-1839.3,-14513.,-16395.
862.0000000000,-5410.1,-4843.7,-1843.9,-14513.,-16395.
863.0000000000,-5415.5,-4846.0,-1846.3,-14512.,-16395.
864.0000000000,-5416.8,-4844.0,-1845.7,-14512.,-16394.
865.0000000000,-5415.9,-4841.0,-1844.2,-14512.,-16394.
866.0000000000,-5417.2,-4842.0,-1845.1,-14512.,-16394.
867.0000000000,-5422.3,-4846.6,-1848.5,-14512.,-16393.
868.0000000000,-5421.4,-4842.5,-1846.3,-14512.,-16393.
869.0000000000,-5418.7,-4838.5,-1843.9,-14511.,-16393.
870.0000000000,-5415.4,-4835.1,-1841.7,-14511.,-16392.
871.0000000000,-5415.1,-4835.8,-1842.2,-14511.,-16392.
872.0000000000,-5413.2,-4833.7,-1841.0,-14511.,-16392.
873.0000000000,-5410.5,-4831.0,-1839.4,-14511.,-16391.
874.0000000000,-5409.2,-4830.5,-1839.1,-14510.,-16391.
875.0000000000,-5406.7,-4828.1,-1837.8,-14510.,-16391.
876.0000000000,-5404.4,-4826.5,-1836.9,-14510.,-16390.
877.0000000000,-5401.5,-4824.1,-1835.5,-14510.,-16390.
878.0000000000,-5398.3,-4821.9,-1834.2,-14510.,-16390.
879.0000000000,-5403.2,-4829.2,-1839.1,-14509.,-16390.
880.0000000000,-5402.7,-4826.6,-1838.0,-14509.,-16389.
881.0000000000,-5406.4,-4830.7,-1841.0,-14509.,-16389.
882.0000000000,-5405.2,-4827.3,-1839.3,-14509.,-16389.
883.0000000000,-5402.4,-4823.9,-1837.3,-14509.,-16388.
884.0000000000,-5399.1,-4821.0,-1835.5,-14508.,-16388.
885.0000000000,-5395.8,-4818.4,-1833.9,-14508.,-16388.
886.0000000000,-5392.5,-4816.2,-1832.5,-14508.,-16387.
887.0000000000,-5389.2,-4814.1,-1831.2,-14508.,-16387.
888.0000000000,-5386.0,-4812.1,-1830.1,-14508.,-16387.
889.0000000000,-5382.9,-4810.3,-1829.0,-14508.,-16386.
890.0000000000,-5379.8,-4808.5,-1828.0,-14507.,-16386.
891.0000000000,-5376.7,-4806.8,-1827.1,-14507.,-16386.
892.0000000000,-5373.7,-4805.2,-1826.2,-14507.,-16385.
893.0000000000,-5370.8,-4803.5,-1825.4,-14507.,-16385.
894.0000000000,-5368.5,-4802.7,-1825.1,-14507.,-16385.
895.0000000000,-5371.1,-4807.2,-1828.4,-14506.,-16384.
896.0000000000,-5370.4,-4805.8,-1828.0,-14506.,-16384.
897.0000000000,-5370.6,-4806.2,-1828.6,-14506.,-16384.
898.0000000000,-5369.5,-4804.9,-1828.2,-14506.,-16383.
899.0000000000,-5367.1,-4802.5,-1826.9,-14506.,-16383.
900.0000000000,-5364.3,-4800.3,-1825.7,-14505.,-16383.
901.0000000000,-5363.7,-4801.0,-1826.4,-14505.,-16382.
902.0000000000,-5361.6,-4799.1,-1825.4,-14505.,-16382.
903.0000000000,-5358.9,-4796.9,-1824.2,-14505.,-16382.
904.0000000000,-5356.5,-4795.6,-1823.5,-14505.,-16381.
905.0000000000,-5353.7,-4793.7,-1822.5,-14505.,-16381.
906.0000000000,-5350.8,-4791.8,-1821.5,-14504.,-16381.
907.0000000000,-5347.8,-4790.1,-1820.6,-14504.,-16381.
908.0000000000,-5348.0,-4792.0,-1822.1,-14504.,-16380.
909.0000000000,-5348.9,-4793.4,-1823.4,-14504.,-16380.
910.0000000000,-5347.3,-4791.2,-1822.4,-14504.,-16380.
911.0000000000,-5344.6,-4788.9,-1821.2,-14503.,-16379.
912.0000000000,-5342.5,-4787.6,-1820.6,-14503.,-16379.
913.0000000000,-5339.7,-4785.7,-1819.5,-14503.,-16379.
914.0000000000,-5336.8,-4783.8,-1818.5,-14503.,-16378.
915.0000000000,-5333.9,-4782.0,-1817.5,-14503.,-16378.
916.0000000000,-5331.0,-4780.4,-1816.6,-14502.,-16378.
917.0000000000,-5328.1,-4778.8,-1815.8,-14502.,-16377.
918.0000000000,-5325.3,-4777.3,-1815.1,-14502.,-16377.
919.0000000000,-5325.7,-4779.5,-1816.8,-14502.,-16377.
920.0000000000,-5323.9,-4777.7,-1816.0,-14502.,-16376.
921.0000000000,-5321.4,-4775.7,-1815.1,-14501.,-16376.
922.0000000000,-5318.6,-4774.0,-1814.2,-14501.,-16376.
923.0000000000,-5315.8,-4772.3,-1813.3,-14501.,-16375.
924.0000000000,-5313.0,-4770.7,-1812.5,-14501.,-16375.
925.0000000000,-5310.3,-4769.2,-1811.8,-14501.,-16375.
926.0000000000,-5307.5,-4767.8,-1811.1,-14500.,-16374.
927.0000000000,-5304.8,-4766.3,-1810.4,-14500.,-16374.
928.0000000000,-5302.1,-4764.9,-1809.8,-14500.,-16374.
929.0000000000,-5299.5,-4763.6,-1809.1,-14500.,-16373.
930.0000000000,-5296.8,-4762.2,-1808.5,-14500.,-16373.
931.0000000000,-5294.2,-4760.9,-1808.0,-14500.,-16373.
932.0000000000,-5291.6,-4759.6,-1807.4,-14499.,-16372.
933.0000000000,-5289.0,-4758.3,-1806.8,-14499.,-16372.
934.0000000000,-5286.5,-4757.0,-1806.3,-14499.,-16372.
935.0000000000,-5283.9,-4755.7,-1805.7,-14499.,-16372.
936.0000000000,-5281.4,-4754.4,-1805.2,-14499.,-16371.
937.0000000000,-5278.9,-4753.1,-1804.7,-14498.,-16371.
938.0000000000,-5276.4,-4751.9,-1804.1,-14498.,-16371.
939.0000000000,-5273.9,-4750.6,-1803.6,-14498.,-16370.
940.0000000000,-5271.4,-4749.4,-1803.1,-14498.,-16370.
941.0000000000,-5269.0,-4748.2,-1802.6,-14498.,-16370.
942.0000000000,-5266.5,-4746.9,-1802.1,-14497.,-16369.
943.0000000000,-5265.0,-4746.7,-1802.3,-14497.,-16369.
944.0000000000,-5263.7,-4746.5,-1802.5,-14497.,-16369.
945.0000000000,-5261.6,-4745.0,-1801.9,-14497.,-16368.
946.0000000000,-5259.3,-4743.5,-1801.3,-14497.,-16368.
947.0000000000,-5256.9,-4742.1,-1800.7,-14496.,-16368.
948.0000000000,-5254.4,-4740.8,-1800.1,-14496.,-16367.
949.0000000000,-5252.0,-4739.5,-1799.6,-14496.,-16367.
950.0000000000,-5249.6,-4738.2,-1799.0,-14496.,-16367.
951.0000000000,-5247.2,-4737.0,-1798.5,-14496.,-16366.
952.0000000000,-5244.8,-4735.8,-1798.0,-14496.,-16366.
953.0000000000,-5242.5,-4734.5,-1797.5,-14495.,-16366.
954.0000000000,-5240.1,-4733.3,-1797.0,-14495.,-16365.
955.0000000000,-5238.7,-4733.2,-1797.2,-14495.,-16365.
956.0000000000,-5237.3,-4732.7,-1797.2,-14495.,-16365.
957.0000000000,-5236.6,-4732.8,-1797.7,-14495.,-16364.
958.0000000000,-5236.7,-4733.6,-1798.6,-14494.,-16364.
959.0000000000,-5235.0,-4731.8,-1797.8,-14494.,-16364.
960.0000000000,-5232.8,-4730.0,-1797.0,-14494.,-16364.
961.0000000000,-5230.5,-4728.4,-1796.2,-14494.,-16363.
962.0000000000,-5230.7,-4730.1,-1797.6,-14494.,-16363.
963.0000000000,-5230.3,-4729.8,-1797.8,-14493.,-16363.
964.0000000000,-5228.5,-4727.9,-1796.9,-14493.,-16362.
965.0000000000,-5226.2,-4726.1,-1796.0,-14493.,-16362.
966.0000000000,-5223.8,-4724.4,-1795.1,-14493.,-16362.
967.0000000000,-5221.4,-4722.9,-1794.4,-14493.,-16361.
968.0000000000,-5219.4,-4722.1,-1794.0,-14492.,-16361.
969.0000000000,-5217.9,-4721.4,-1793.9,-14492.,-16361.
970.0000000000,-5215.7,-4720.0,-1793.2,-14492.,-16360.
971.0000000000,-5213.4,-4718.5,-1792.5,-14492.,-16360.
972.0000000000,-5211.1,-4717.1,-1791.8,-14492.,-16360.
973.0000000000,-5209.1,-4716.2,-1791.5,-14491.,-16359.
974.0000000000,-5206.9,-4714.9,-1790.9,-14491.,-16359.
975.0000000000,-5204.6,-4713.6,-1790.3,-14491.,-16359.
976.0000000000,-5202.3,-4712.3,-1789.7,-14491.,-16358.
977.0000000000,-5200.0,-4711.1,-1789.2,-14491.,-16358.
978.0000000000,-5197.8,-4709.9,-1788.6,-14490.,-16358.
979.0000000000,-5195.5,-4708.7,-1788.1,-14490.,-16357.
980.0000000000,-5193.3,-4707.5,-1787.6,-14490.,-16357.
981.0000000000,-5191.1,-4706.4,-1787.1,-14490.,-16357.
982.0000000000,-5188.9,-4705.2,-1786.6,-14490.,-16357.
983.0000000000,-5188.2,-4705.9,-1787.4,-14490.,-16356.
984.0000000000,-5186.5,-4704.6,-1786.9,-14489.,-16356.
985.0000000000,-5185.3,-4704.2,-1787.0,-14489.,-16356.
986.0000000000,-5183.4,-4702.8,-1786.4,-14489.,-16355.
987.0000000000,-5181.3,-4701.4,-1785.7,-14489.,-16355.
988.0000000000,-5179.1,-4700.1,-1785.1,-14489.,-16355.
989.0000000000,-5176.9,-4698.9,-1784.6,-14488.,-16354.
990.0000000000,-5174.7,-4697.6,-1784.0,-14488.,-16354.
991.0000000000,-5172.5,-4696.5,-1783.5,-14488.,-16354.
992.0000000000,-5170.3,-4695.3,-1783.0,-14488.,-16353.
993.0000000000,-5168.2,-4694.1,-1782.5,-14488.,-16353.
994.0000000000,-5166.0,-4693.0,-1782.0,-14487.,-16353.
995.0000000000,-5163.9,-4691.9,-1781.6,-14487.,-16352.
996.0000000000,-5161.8,-4690.8,-1781.1,-14487.,-16352.
997.0000000000,-5159.7,-4689.7,-1780.7,-14487.,-16352.
998.0000000000,-5157.6,-4688.6,-1780.2,-14487.,-16351.
999.0000000000,-5155.5,-4687.5,-1779.8,-14486.,-16351.
1000.000000000,-5154.1,-4687.1,-1779.8,-14486.,-16351.
1001.000000000,-5152.2,-4686.0,-1779.4,-14486.,-16350.
1002.000000000,-5150.2,-4684.8,-1778.9,-14486.,-16350.
1003.000000000,-5148.1,-4683.7,-1778.4,-14486.,-16350.
1004.000000000,-5146.1,-4682.5,-1778.0,-14485.,-16350.
1005.000000000,-5144.0,-4681.4,-1777.5,-14485.,-16349.
1006.000000000,-5142.0,-4680.4,-1777.1,-14485.,-16349.
1007.000000000,-5139.9,-4679.3,-1776.7,-14485.,-16349.
1008.000000000,-5137.9,-4678.2,-1776.2,-14485.,-16348.
1009.000000000,-5135.9,-4677.2,-1775.8,-14485.,-16348.
1010.000000000,-5133.9,-4676.1,-1775.4,-14484.,-16348.
1011.000000000,-5131.9,-4675.1,-1775.0,-14484.,-16347.
1012.000000000,-5137.2,-4682.5,-1780.2,-14484.,-16347.
1013.000000000,-5138.5,-4682.0,-1780.5,-14484.,-16347.
1014.000000000,-5137.3,-4679.7,-1779.5,-14484.,-16346.
1015.000000000,-5135.4,-4677.6,-1778.4,-14483.,-16346.
1016.000000000,-5133.2,-4675.8,-1777.4,-14483.,-16346.
1017.000000000,-5131.0,-4674.2,-1776.5,-14483.,-16345.
1018.000000000,-5128.7,-4672.8,-1775.7,-14483.,-16345.
1019.000000000,-5126.6,-4671.4,-1775.0,-14483.,-16345.
1020.000000000,-5124.4,-4670.1,-1774.4,-14482.,-16345.
1021.000000000,-5122.3,-4668.9,-1773.8,-14482.,-16344.
1022.000000000,-5120.2,-4667.7,-1773.2,-14482.,-16344.
1023.000000000,-5118.1,-4666.5,-1772.6,-14482.,-16344.
1024.000000000,-5116.0,-4665.4,-1772.1,-14482.,-16343.
1025.000000000,-5114.4,-4664.8,-1771.9,-14481.,-16343.
1026.000000000,-5113.3,-4664.6,-1772.1,-14481.,-16343.
1027.000000000,-5126.6,-4680.9,-1783.1,-14481.,-16342.
1028.000000000,-5135.7,-4685.9,-1787.4,-14481.,-16342.
1029.000000000,-5136.7,-4681.5,-1785.4,-14481.,-16342.
1030.000000000,-5135.0,-4677.5,-1783.0,-14480.,-16341.
1031.000000000,-5132.5,-4674.2,-1781.0,-14480.,-16341.
1032.000000000,-5129.8,-4671.6,-1779.2,-14480.,-16341.
1033.000000000,-5127.7,-4670.1,-1778.2,-14480.,-16340.
1034.000000000,-5134.0,-4678.4,-1783.6,-14480.,-16340.
1035.000000000,-5134.1,-4675.6,-1782.3,-14479.,-16340.
1036.000000000,-5132.2,-4672.5,-1780.4,-14479.,-16339.
1037.000000000,-5129.7,-4669.8,-1778.7,-14479.,-16339.
1038.000000000,-5127.1,-4667.6,-1777.2,-14479.,-16339.
1039.000000000,-5124.4,-4665.7,-1776.0,-14479.,-16339.
1040.000000000,-5121.8,-4663.9,-1774.8,-14479.,-16338.
1041.000000000,-5119.7,-4662.7,-1774.1,-14478.,-16338.
1042.000000000,-5117.6,-4661.6,-1773.4,-14478.,-16338.
1043.000000000,-5115.3,-4660.0,-1772.5,-14478.,-16337.
1044.000000000,-5113.0,-4658.6,-1771.6,-14478.,-16337.
1045.000000000,-5110.6,-4657.2,-1770.8,-14478.,-16337.
1046.000000000,-5108.2,-4655.9,-1770.1,-14477.,-16336.
1047.000000000,-5105.9,-4654.6,-1769.4,-14477.,-16336.
1048.000000000,-5103.8,-4653.6,-1768.9,-14477.,-16336.
1049.000000000,-5102.2,-4653.1,-1768.7,-14477.,-16335.
1050.000000000,-5100.3,-4652.0,-1768.2,-14477.,-16335.
1051.000000000,-5098.4,-4651.0,-1767.7,-14476.,-16335.
1052.000000000,-5096.2,-4649.7,-1767.1,-14476.,-16334.
1053.000000000,-5094.0,-4648.5,-1766.5,-14476.,-16334.
1054.000000000,-5091.8,-4647.3,-1765.9,-14476.,-16334.
1055.000000000,-5089.6,-4646.2,-1765.3,-14476.,-16334.
1056.000000000,-5087.4,-4645.1,-1764.8,-14475.,-16333.
1057.000000000,-5085.3,-4644.0,-1764.2,-14475.,-16333.
1058.000000000,-5083.1,-4642.9,-1763.7,-14475.,-16333.
1059.000000000,-5081.0,-4641.8,-1763.2,-14475.,-16332.
1060.000000000,-5079.2,-4641.1,-1763.0,-14475.,-16332.
1061.000000000,-5078.4,-4641.5,-1763.5,-14474.,-16332.
1062.000000000,-5082.2,-4646.7,-1767.2,-14474.,-16331.
1063.000000000,-5082.1,-4645.2,-1766.7,-14474.,-16331.
1064.000000000,-5080.4,-4643.0,-1765.6,-14474.,-16331.
1065.000000000,-5078.3,-4641.2,-1764.6,-14474.,-16330.
1066.000000000,-5076.0,-4639.6,-1763.7,-14473.,-16330.
1067.000000000,-5073.8,-4638.2,-1762.9,-14473.,-16330.
1068.000000000,-5071.5,-4636.9,-1762.2,-14473.,-16330.
1069.000000000,-5069.3,-4635.6,-1761.5,-14473.,-16329.
1070.000000000,-5067.1,-4634.4,-1760.9,-14473.,-16329.
1071.000000000,-5065.0,-4633.3,-1760.3,-14472.,-16329.
1072.000000000,-5062.8,-4632.1,-1759.8,-14472.,-16328.
1073.000000000,-5060.7,-4631.1,-1759.2,-14472.,-16328.
1074.000000000,-5058.6,-4630.0,-1758.7,-14472.,-16328.
1075.000000000,-5056.6,-4628.9,-1758.2,-14472.,-16327.
1076.000000000,-5054.5,-4627.9,-1757.8,-14472.,-16327.
1077.000000000,-5058.8,-4634.3,-1762.2,-14471.,-16327.
1078.000000000,-5058.7,-4632.7,-1761.7,-14471.,-16326.
1079.000000000,-5057.1,-4630.6,-1760.6,-14471.,-16326.
1080.000000000,-5055.1,-4628.9,-1759.7,-14471.,-16326.
1081.000000000,-5052.9,-4627.3,-1758.8,-14471.,-16325.
1082.000000000,-5050.7,-4625.9,-1758.1,-14470.,-16325.
1083.000000000,-5048.5,-4624.7,-1757.4,-14470.,-16325.
1084.000000000,-5046.4,-4623.5,-1756.7,-14470.,-16325.
1085.000000000,-5044.3,-4622.3,-1756.1,-14470.,-16324.
1086.000000000,-5042.2,-4621.2,-1755.6,-14470.,-16324.
1087.000000000,-5040.1,-4620.1,-1755.0,-14469.,-16324.
1088.000000000,-5038.1,-4619.0,-1754.5,-14469.,-16323.
1089.000000000,-5036.1,-4618.0,-1754.0,-14469.,-16323.
1090.000000000,-5034.1,-4617.0,-1753.6,-14469.,-16323.
1091.000000000,-5037.4,-4622.3,-1757.3,-14469.,-16322.
1092.000000000,-5038.2,-4622.1,-1757.6,-14468.,-16322.
1093.000000000,-5036.9,-4620.1,-1756.7,-14468.,-16322.
1094.000000000,-5035.0,-4618.3,-1755.7,-14468.,-16321.
1095.000000000,-5032.9,-4616.7,-1754.8,-14468.,-16321.
1096.000000000,-5030.7,-4615.3,-1754.0,-14468.,-16321.
1097.000000000,-5028.7,-4614.1,-1753.4,-14467.,-16321.
1098.000000000,-5027.6,-4614.0,-1753.5,-14467.,-16320.
1099.000000000,-5025.8,-4612.8,-1752.9,-14467.,-16320.
1100.000000000,-5023.8,-4611.5,-1752.2,-14467.,-16320.
1101.000000000,-5021.8,-4610.3,-1751.6,-14467.,-16319.
1102.000000000,-5019.8,-4609.2,-1751.0,-14466.,-16319.
1103.000000000,-5017.8,-4608.1,-1750.5,-14466.,-16319.
1104.000000000,-5015.8,-4607.0,-1750.0,-14466.,-16318.
1105.000000000,-5013.8,-4606.0,-1749.5,-14466.,-16318.
1106.000000000,-5011.8,-4605.0,-1749.0,-14466.,-16318.
1107.000000000,-5009.9,-4604.0,-1748.5,-14465.,-16317.
1108.000000000,-5008.0,-4603.0,-1748.1,-14465.,-16317.
1109.000000000,-5006.0,-4602.1,-1747.7,-14465.,-16317.
1110.000000000,-5004.1,-4601.1,-1747.2,-14465.,-16317.
1111.000000000,-5002.2,-4600.2,-1746.8,-14465.,-16316.
1112.000000000,-5000.4,-4599.2,-1746.4,-14465.,-16316.
1113.000000000,-4998.5,-4598.3,-1746.0,-14464.,-16316.
1114.000000000,-4996.6,-4597.4,-1745.6,-14464.,-16315.
1115.000000000,-4994.8,-4596.5,-1745.2,-14464.,-16315.
1116.000000000,-4993.0,-4595.5,-1744.9,-14464.,-16315.
1117.000000000,-4991.1,-4594.6,-1744.5,-14464.,-16314.
1118.000000000,-4989.3,-4593.7,-1744.1,-14463.,-16314.
1119.000000000,-4987.5,-4592.8,-1743.7,-14463.,-16314.
1120.000000000,-4985.7,-4591.9,-1743.4,-14463.,-16313.
1121.000000000,-4983.9,-4591.0,-1743.0,-14463.,-16313.
1122.000000000,-4985.4,-4594.0,-1745.2,-14463.,-16313.
1123.000000000,-4984.6,-4592.8,-1744.8,-14462.,-16313.
1124.000000000,-4983.0,-4591.4,-1744.1,-14462.,-16312.
1125.000000000,-4981.3,-4590.1,-1743.5,-14462.,-16312.
1126.000000000,-4979.4,-4588.9,-1742.9,-14462.,-16312.
1127.000000000,-4977.6,-4587.9,-1742.4,-14462.,-16311.
1128.000000000,-4975.7,-4586.8,-1741.9,-14461.,-16311.
1129.000000000,-4973.9,-4585.8,-1741.4,-14461.,-16311.
1130.000000000,-4972.1,-4584.9,-1741.0,-14461.,-16310.
1131.000000000,-4970.3,-4583.9,-1740.6,-14461.,-16310.
1132.000000000,-4968.5,-4583.0,-1740.2,-14461.,-16310.
1133.000000000,-4966.7,-4582.1,-1739.8,-14460.,-16309.
1134.000000000,-4965.0,-4581.2,-1739.4,-14460.,-16309.
1135.000000000,-4963.2,-4580.3,-1739.0,-14460.,-16309.
1136.000000000,-4961.5,-4579.4,-1738.6,-14460.,-16309.
1137.000000000,-4959.8,-4578.5,-1738.3,-14460.,-16308.
1138.000000000,-4958.1,-4577.6,-1737.9,-14459.,-16308.
1139.000000000,-4956.4,-4576.8,-1737.5,-14459.,-16308.
1140.000000000,-4954.7,-4575.9,-1737.2,-14459.,-16307.
1141.000000000,-4953.0,-4575.0,-1736.8,-14459.,-16307.
1142.000000000,-4951.3,-4574.2,-1736.5,-14459.,-16307.
1143.000000000,-4949.6,-4573.3,-1736.1,-14458.,-16306.
1144.000000000,-4947.9,-4572.5,-1735.8,-14458.,-16306.
1145.000000000,-4946.3,-4571.6,-1735.5,-14458.,-16306.
1146.000000000,-4944.6,-4570.8,-1735.1,-14458.,-16306.
1147.000000000,-4943.0,-4570.0,-1734.8,-14458.,-16305.
1148.000000000,-4942.6,-4570.6,-1735.4,-14457.,-16305.
1149.000000000,-4944.8,-4573.7,-1737.8,-14457.,-16305.
1150.000000000,-4944.3,-4572.3,-1737.3,-14457.,-16304.
1151.000000000,-4942.9,-4570.7,-1736.5,-14457.,-16304.
1152.000000000,-4941.2,-4569.4,-1735.8,-14457.,-16304.
1153.000000000,-4939.4,-4568.2,-1735.2,-14457.,-16303.
1154.000000000,-4937.7,-4567.1,-1734.6,-14456.,-16303.
1155.000000000,-4935.9,-4566.0,-1734.1,-14456.,-16303.
1156.000000000,-4934.2,-4565.0,-1733.6,-14456.,-16302.
1157.000000000,-4932.5,-4564.1,-1733.2,-14456.,-16302.
1158.000000000,-4930.8,-4563.2,-1732.7,-14456.,-16302.
1159.000000000,-4929.1,-4562.3,-1732.3,-14455.,-16302.
1160.000000000,-4927.5,-4561.4,-1731.9,-14455.,-16301.
1161.000000000,-4925.8,-4560.5,-1731.5,-14455.,-16301.
1162.000000000,-4924.2,-4559.6,-1731.2,-14455.,-16301.
1163.000000000,-4928.3,-4565.5,-1735.2,-14455.,-16300.
1164.000000000,-4932.0,-4568.4,-1737.6,-14454.,-16300.
1165.000000000,-4937.3,-4572.7,-1740.9,-14454.,-16300.
1166.000000000,-4943.0,-4576.3,-1743.9,-14454.,-16299.
1167.000000000,-4946.4,-4577.0,-1744.8,-14454.,-16299.
1168.000000000,-4945.9,-4573.6,-1742.9,-14454.,-16299.
1169.000000000,-4944.0,-4570.6,-1741.0,-14453.,-16299.
1170.000000000,-4941.8,-4568.1,-1739.4,-14453.,-16298.
1171.000000000,-4939.5,-4566.1,-1738.0,-14453.,-16298.
1172.000000000,-4937.4,-4564.4,-1736.8,-14453.,-16298.
1173.000000000,-4935.3,-4562.9,-1735.8,-14453.,-16297.
1174.000000000,-4935.8,-4564.6,-1736.9,-14452.,-16297.
1175.000000000,-4934.6,-4563.0,-1736.0,-14452.,-16297.
1176.000000000,-4932.7,-4561.3,-1734.9,-14452.,-16296.
1177.000000000,-4930.7,-4559.8,-1734.0,-14452.,-16296.
1178.000000000,-4928.7,-4558.5,-1733.2,-14452.,-16296.
1179.000000000,-4927.1,-4557.6,-1732.7,-14451.,-16296.
1180.000000000,-4925.2,-4556.4,-1732.0,-14451.,-16295.
1181.000000000,-4923.3,-4555.3,-1731.3,-14451.,-16295.
1182.000000000,-4921.4,-4554.2,-1730.7,-14451.,-16295.
1183.000000000,-4919.5,-4553.1,-1730.1,-14451.,-16294.
1184.000000000,-4917.6,-4552.1,-1729.5,-14450.,-16294.
1185.000000000,-4915.8,-4551.1,-1729.0,-14450.,-16294.
1186.000000000,-4914.0,-4550.1,-1728.5,-14450.,-16293.
1187.000000000,-4912.2,-4549.3,-1728.1,-14450.,-16293.
1188.000000000,-4910.4,-4548.4,-1727.6,-14450.,-16293.
1189.000000000,-4908.6,-4547.4,-1727.1,-14449.,-16293.
1190.000000000,-4906.9,-4546.5,-1726.7,-14449.,-16292.
1191.000000000,-4905.1,-4545.7,-1726.3,-14449.,-16292.
1192.000000000,-4903.3,-4544.8,-1725.9,-14449.,-16292.
1193.000000000,-4901.6,-4543.9,-1725.5,-14449.,-16291.
1194.000000000,-4899.9,-4543.1,-1725.1,-14449.,-16291.
1195.000000000,-4898.2,-4542.2,-1724.7,-14448.,-16291.
1196.000000000,-4896.5,-4541.4,-1724.3,-14448.,-16290.
1197.000000000,-4894.9,-4540.7,-1724.0,-14448.,-16290.
1198.000000000,-4893.2,-4539.8,-1723.6,-14448.,-16290.
1199.000000000,-4893.9,-4541.8,-1725.1,-14448.,-16289.
1200.000000000,-4892.9,-4540.7,-1724.7,-14447.,-16289.
1201.000000000,-4891.4,-4539.5,-1724.1,-14447.,-16289.
1202.000000000,-4889.8,-4538.4,-1723.6,-14447.,-16289.
1203.000000000,-4903.7,-4555.9,-1735.3,-14447.,-16288.
1204.000000000,-4910.2,-4557.5,-1737.3,-14447.,-16288.
1205.000000000,-4910.7,-4553.7,-1735.4,-14446.,-16288.
1206.000000000,-4909.2,-4550.4,-1733.4,-14446.,-16287.
1207.000000000,-4907.1,-4547.7,-1731.7,-14446.,-16287.
1208.000000000,-4904.9,-4545.6,-1730.2,-14446.,-16287.
1209.000000000,-4902.7,-4543.8,-1728.9,-14446.,-16287.
1210.000000000,-4900.8,-4542.4,-1728.0,-14445.,-16286.
1211.000000000,-4898.7,-4541.0,-1727.0,-14445.,-16286.
1212.000000000,-4896.6,-4539.6,-1726.1,-14445.,-16286.
1213.000000000,-4896.2,-4540.1,-1726.5,-14445.,-16285.
1214.000000000,-4894.6,-4538.8,-1725.7,-14445.,-16285.
1215.000000000,-4892.8,-4537.4,-1724.9,-14444.,-16285.
1216.000000000,-4890.9,-4536.2,-1724.1,-14444.,-16284.
1217.000000000,-4889.0,-4535.1,-1723.4,-14444.,-16284.
1218.000000000,-4887.1,-4534.0,-1722.8,-14444.,-16284.
1219.000000000,-4885.3,-4533.0,-1722.2,-14444.,-16284.
1220.000000000,-4883.4,-4532.0,-1721.7,-14443.,-16283.
1221.000000000,-4881.5,-4531.0,-1721.1,-14443.,-16283.
1222.000000000,-4879.7,-4530.0,-1720.6,-14443.,-16283.
1223.000000000,-4877.9,-4529.1,-1720.1,-14443.,-16282.
1224.000000000,-4876.1,-4528.2,-1719.7,-14443.,-16282.
1225.000000000,-4874.8,-4527.9,-1719.6,-14442.,-16282.
1226.000000000,-4873.2,-4527.0,-1719.2,-14442.,-16281.
1227.000000000,-4871.5,-4526.1,-1718.7,-14442.,-16281.
1228.000000000,-4869.8,-4525.2,-1718.3,-14442.,-16281.
1229.000000000,-4868.1,-4524.4,-1717.9,-14442.,-16281.
1230.000000000,-4866.4,-4523.5,-1717.5,-14441.,-16280.
1231.000000000,-4865.5,-4523.6,-1717.7,-14441.,-16280.
1232.000000000,-4864.6,-4523.3,-1717.7,-14441.,-16280.
1233.000000000,-4863.1,-4522.3,-1717.2,-14441.,-16279.
1234.000000000,-4863.3,-4523.5,-1718.2,-14441.,-16279.
1235.000000000,-4867.2,-4528.3,-1721.6,-14440.,-16279.
1236.000000000,-4868.1,-4527.7,-1721.7,-14440.,-16278.
1237.000000000,-4867.0,-4525.7,-1720.6,-14440.,-16278.
1238.000000000,-4865.3,-4523.9,-1719.6,-14440.,-16278.
1239.000000000,-4863.4,-4522.4,-1718.7,-14440.,-16278.
1240.000000000,-4861.5,-4521.1,-1717.9,-14440.,-16277.
1241.000000000,-4859.6,-4519.9,-1717.2,-14439.,-16277.
1242.000000000,-4857.8,-4518.8,-1716.5,-14439.,-16277.
1243.000000000,-4856.0,-4517.8,-1716.0,-14439.,-16276.
1244.000000000,-4854.2,-4516.8,-1715.4,-14439.,-16276.
1245.000000000,-4852.5,-4515.9,-1714.9,-14439.,-16276.
1246.000000000,-4851.0,-4515.2,-1714.6,-14438.,-16275.
1247.000000000,-4849.3,-4514.3,-1714.1,-14438.,-16275.
1248.000000000,-4848.2,-4514.1,-1714.1,-14438.,-16275.
1249.000000000,-4856.8,-4525.2,-1721.5,-14438.,-16275.
1250.000000000,-4860.5,-4525.8,-1722.7,-14438.,-16274.
1251.000000000,-4860.3,-4523.3,-1721.4,-14437.,-16274.
1252.000000000,-4858.8,-4520.8,-1719.9,-14437.,-16274.
1253.000000000,-4856.8,-4518.7,-1718.6,-14437.,-16273.
1254.000000000,-4854.8,-4517.0,-1717.5,-14437.,-16273.
1255.000000000,-4852.8,-4515.5,-1716.5,-14437.,-16273.
1256.000000000,-4850.8,-4514.2,-1715.7,-14436.,-16273.
1257.000000000,-4848.8,-4513.0,-1714.9,-14436.,-16272.
1258.000000000,-4846.9,-4511.9,-1714.2,-14436.,-16272.
1259.000000000,-4845.0,-4510.8,-1713.5,-14436.,-16272.
1260.000000000,-4843.3,-4509.9,-1713.0,-14436.,-16271.
1261.000000000,-4841.5,-4509.0,-1712.5,-14435.,-16271.
1262.000000000,-4839.8,-4508.0,-1711.9,-14435.,-16271.
1263.000000000,-4838.0,-4507.1,-1711.4,-14435.,-16270.
1264.000000000,-4836.3,-4506.2,-1711.0,-14435.,-16270.
1265.000000000,-4834.5,-4505.3,-1710.5,-14435.,-16270.
1266.000000000,-4832.8,-4504.5,-1710.1,-14434.,-16270.
1267.000000000,-4833.4,-4506.3,-1711.4,-14434.,-16269.
1268.000000000,-4832.4,-4505.3,-1711.0,-14434.,-16269.
1269.000000000,-4830.8,-4504.1,-1710.4,-14434.,-16269.
1270.000000000,-4829.2,-4503.0,-1709.8,-14434.,-16268.
1271.000000000,-4827.5,-4502.0,-1709.3,-14433.,-16268.
1272.000000000,-4825.8,-4501.1,-1708.8,-14433.,-16268.
1273.000000000,-4826.2,-4502.8,-1710.0,-14433.,-16268.
1274.000000000,-4842.1,-4521.8,-1722.8,-14433.,-16267.
1275.000000000,-4846.4,-4519.6,-1722.4,-14433.,-16267.
1276.000000000,-4846.2,-4515.8,-1720.4,-14432.,-16267.
1277.000000000,-4844.5,-4512.6,-1718.4,-14432.,-16266.
1278.000000000,-4842.3,-4510.1,-1716.7,-14432.,-16266.
1279.000000000,-4840.1,-4508.1,-1715.2,-14432.,-16266.
1280.000000000,-4837.9,-4506.3,-1714.0,-14432.,-16265.
1281.000000000,-4835.7,-4504.8,-1712.9,-14432.,-16265.
1282.000000000,-4833.6,-4503.4,-1711.9,-14431.,-16265.
1283.000000000,-4831.6,-4502.2,-1711.1,-14431.,-16265.
1284.000000000,-4829.6,-4501.0,-1710.3,-14431.,-16264.
1285.000000000,-4827.7,-4499.9,-1709.6,-14431.,-16264.
1286.000000000,-4825.8,-4498.8,-1709.0,-14431.,-16264.
1287.000000000,-4823.9,-4497.9,-1708.4,-14430.,-16263.
1288.000000000,-4822.1,-4496.9,-1707.8,-14430.,-16263.
1289.000000000,-4820.3,-4496.0,-1707.3,-14430.,-16263.
1290.000000000,-4818.5,-4495.1,-1706.8,-14430.,-16263.
1291.000000000,-4816.7,-4494.2,-1706.3,-14430.,-16262.
1292.000000000,-4815.0,-4493.3,-1705.8,-14429.,-16262.
1293.000000000,-4813.2,-4492.5,-1705.4,-14429.,-16262.
1294.000000000,-4811.5,-4491.6,-1704.9,-14429.,-16261.
1295.000000000,-4809.8,-4490.8,-1704.5,-14429.,-16261.
1296.000000000,-4808.1,-4490.0,-1704.1,-14429.,-16261.
1297.000000000,-4806.4,-4489.2,-1703.7,-14428.,-16260.
1298.000000000,-4804.7,-4488.4,-1703.4,-14428.,-16260.
1299.000000000,-4803.1,-4487.7,-1703.0,-14428.,-16260.
1300.000000000,-4801.4,-4486.9,-1702.6,-14428.,-16260.
1301.000000000,-4799.8,-4486.1,-1702.3,-14428.,-16259.
1302.000000000,-4798.2,-4485.4,-1701.9,-14427.,-16259.
1303.000000000,-4796.6,-4484.7,-1701.6,-14427.,-16259.
1304.000000000,-4796.8,-4486.0,-1702.6,-14427.,-16258.
1305.000000000,-4795.9,-4485.3,-1702.4,-14427.,-16258.
1306.000000000,-4794.5,-4484.2,-1701.9,-14427.,-16258.
1307.000000000,-4793.0,-4483.3,-1701.5,-14426.,-16258.
1308.000000000,-4791.4,-4482.4,-1701.0,-14426.,-16257.
1309.000000000,-4789.7,-4481.6,-1700.6,-14426.,-16257.
1310.000000000,-4788.1,-4480.7,-1700.2,-14426.,-16257.
1311.000000000,-4786.5,-4479.9,-1699.8,-14426.,-16256.
1312.000000000,-4785.0,-4479.2,-1699.4,-14425.,-16256.
1313.000000000,-4783.4,-4478.4,-1699.1,-14425.,-16256.
1314.000000000,-4781.8,-4477.6,-1698.7,-14425.,-16256.
1315.000000000,-4780.3,-4476.9,-1698.4,-14425.,-16255.
1316.000000000,-4778.7,-4476.1,-1698.0,-14425.,-16255.
1317.000000000,-4777.2,-4475.4,-1697.7,-14424.,-16255.
1318.000000000,-4775.7,-4474.7,-1697.4,-14424.,-16254.
1319.000000000,-4774.2,-4474.0,-1697.1,-14424.,-16254.
1320.000000000,-4772.7,-4473.3,-1696.8,-14424.,-16254.
1321.000000000,-4777.4,-4479.9,-1701.3,-14424.,-16253.
1322.000000000,-4783.1,-4484.9,-1705.1,-14424.,-16253.
1323.000000000,-4785.7,-4485.1,-1705.7,-14423.,-16253.
1324.000000000,-4785.6,-4483.0,-1704.7,-14423.,-16253.
1325.000000000,-4787.9,-4485.2,-1706.3,-14423.,-16252.
1326.000000000,-4788.4,-4484.3,-1706.0,-14423.,-16252.
1327.000000000,-4787.6,-4482.5,-1705.0,-14423.,-16252.
1328.000000000,-4799.0,-4496.0,-1713.8,-14422.,-16251.
1329.000000000,-4802.6,-4494.8,-1713.7,-14422.,-16251.
1330.000000000,-4804.6,-4493.9,-1713.4,-14422.,-16251.
1331.000000000,-4806.5,-4494.1,-1713.7,-14422.,-16251.
1332.000000000,-4805.4,-4490.9,-1711.6,-14422.,-16250.
1333.000000000,-4803.7,-4488.4,-1709.8,-14421.,-16250.
1334.000000000,-4801.4,-4486.0,-1708.1,-14421.,-16250.
1335.000000000,-4799.1,-4483.9,-1706.5,-14421.,-16249.
1336.000000000,-4797.1,-4482.4,-1705.3,-14421.,-16249.
1337.000000000,-4795.8,-4481.9,-1704.9,-14421.,-16249.
1338.000000000,-4794.4,-4480.8,-1704.1,-14420.,-16249.
1339.000000000,-4793.4,-4480.4,-1703.8,-14420.,-16248.
1340.000000000,-4792.1,-4479.5,-1703.2,-14420.,-16248.
1341.000000000,-4790.8,-4478.6,-1702.6,-14420.,-16248.
1342.000000000,-4790.9,-4479.4,-1703.2,-14420.,-16247.
1343.000000000,-4789.5,-4478.0,-1702.3,-14419.,-16247.
1344.000000000,-4787.7,-4476.4,-1701.3,-14419.,-16247.
1345.000000000,-4785.7,-4475.1,-1700.4,-14419.,-16247.
1346.000000000,-4783.7,-4473.9,-1699.6,-14419.,-16246.
1347.000000000,-4781.8,-4472.8,-1698.9,-14419.,-16246.
1348.000000000,-4779.8,-4471.7,-1698.2,-14418.,-16246.
1349.000000000,-4777.9,-4470.7,-1697.6,-14418.,-16245.
1350.000000000,-4776.7,-4470.6,-1697.6,-14418.,-16245.
1351.000000000,-4775.0,-4469.6,-1697.0,-14418.,-16245.
1352.000000000,-4774.9,-4470.6,-1697.8,-14418.,-16245.
1353.000000000,-4773.8,-4469.7,-1697.3,-14418.,-16244.
1354.000000000,-4772.9,-4469.4,-1697.2,-14417.,-16244.
1355.000000000,-4771.3,-4468.2,-1696.6,-14417.,-16244.
1356.000000000,-4769.6,-4467.1,-1695.9,-14417.,-16243.
1357.000000000,-4767.7,-4466.1,-1695.3,-14417.,-16243.
1358.000000000,-4765.9,-4465.1,-1694.8,-14417.,-16243.
1359.000000000,-4764.1,-4464.2,-1694.2,-14416.,-16243.
1360.000000000,-4762.4,-4463.3,-1693.8,-14416.,-16242.
1361.000000000,-4760.6,-4462.5,-1693.3,-14416.,-16242.
1362.000000000,-4758.9,-4461.7,-1692.9,-14416.,-16242.
1363.000000000,-4757.1,-4460.9,-1692.4,-14416.,-16241.
1364.000000000,-4763.6,-4469.8,-1698.4,-14415.,-16241.
1365.000000000,-4783.1,-4490.5,-1712.6,-14415.,-16241.
1366.000000000,-4789.7,-4488.9,-1712.8,-14415.,-16241.
1367.000000000,-4789.9,-4483.8,-1710.0,-14415.,-16240.
1368.000000000,-4788.0,-4479.7,-1707.3,-14415.,-16240.
1369.000000000,-4785.6,-4476.6,-1705.1,-14414.,-16240.
1370.000000000,-4783.0,-4474.0,-1703.2,-14414.,-16239.
1371.000000000,-4780.5,-4471.9,-1701.6,-14414.,-16239.
1372.000000000,-4778.1,-4470.1,-1700.2,-14414.,-16239.
1373.000000000,-4775.8,-4468.5,-1699.0,-14414.,-16239.
1374.000000000,-4773.5,-4467.1,-1698.0,-14413.,-16238.
1375.000000000,-4771.4,-4465.8,-1697.0,-14413.,-16238.
1376.000000000,-4769.3,-4464.6,-1696.2,-14413.,-16238.
1377.000000000,-4767.2,-4463.5,-1695.4,-14413.,-16237.
1378.000000000,-4765.2,-4462.5,-1694.7,-14413.,-16237.
1379.000000000,-4763.2,-4461.4,-1694.0,-14412.,-16237.
1380.000000000,-4761.3,-4460.5,-1693.4,-14412.,-16237.
1381.000000000,-4759.4,-4459.5,-1692.8,-14412.,-16236.
1382.000000000,-4757.5,-4458.6,-1692.3,-14412.,-16236.
1383.000000000,-4755.6,-4457.7,-1691.8,-14412.,-16236.
1384.000000000,-4753.7,-4456.9,-1691.3,-14412.,-16235.
1385.000000000,-4751.9,-4456.0,-1690.8,-14411.,-16235.
1386.000000000,-4750.1,-4455.2,-1690.4,-14411.,-16235.
1387.000000000,-4748.3,-4454.4,-1689.9,-14411.,-16235.
1388.000000000,-4746.5,-4453.6,-1689.5,-14411.,-16234.
1389.000000000,-4744.7,-4452.9,-1689.1,-14411.,-16234.
1390.000000000,-4743.0,-4452.1,-1688.8,-14410.,-16234.
1391.000000000,-4741.3,-4451.4,-1688.4,-14410.,-16234.
1392.000000000,-4739.6,-4450.6,-1688.0,-14410.,-16233.
1393.000000000,-4737.9,-4449.9,-1687.6,-14410.,-16233.
1394.000000000,-4736.2,-4449.2,-1687.3,-14410.,-16233.
1395.000000000,-4734.5,-4448.4,-1686.9,-14409.,-16232.
1396.000000000,-4732.8,-4447.7,-1686.6,-14409.,-16232.
1397.000000000,-4731.2,-4447.0,-1686.3,-14409.,-16232.
1398.000000000,-4729.5,-4446.3,-1685.9,-14409.,-16232.
1399.000000000,-4727.9,-4445.6,-1685.6,-14409.,-16231.
1400.000000000,-4726.3,-4444.9,-1685.3,-14408.,-16231.
1401.000000000,-4724.7,-4444.2,-1685.0,-14408.,-16231.
1402.000000000,-4723.1,-4443.5,-1684.7,-14408.,-16230.
1403.000000000,-4721.5,-4442.8,-1684.4,-14408.,-16230.
1404.000000000,-4723.5,-4446.4,-1686.9,-14408.,-16230.
1405.000000000,-4723.1,-4445.5,-1686.6,-14407.,-16230.
1406.000000000,-4721.9,-4444.3,-1686.0,-14407.,-16229.
1407.000000000,-4720.8,-4443.7,-1685.8,-14407.,-16229.
1408.000000000,-4719.3,-4442.7,-1685.3,-14407.,-16229.
1409.000000000,-4717.7,-4441.7,-1684.7,-14407.,-16228.
1410.000000000,-4721.4,-4447.2,-1688.4,-14406.,-16228.
1411.000000000,-4721.6,-4445.9,-1688.0,-14406.,-16228.
1412.000000000,-4720.4,-4444.2,-1687.1,-14406.,-16228.
1413.000000000,-4718.8,-4442.8,-1686.3,-14406.,-16227.
1414.000000000,-4717.0,-4441.5,-1685.5,-14406.,-16227.
1415.000000000,-4715.3,-4440.4,-1684.8,-14406.,-16227.
1416.000000000,-4713.6,-4439.4,-1684.2,-14405.,-16226.
1417.000000000,-4711.9,-4438.5,-1683.7,-14405.,-16226.
1418.000000000,-4710.2,-4437.6,-1683.2,-14405.,-16226.
1419.000000000,-4708.6,-4436.8,-1682.8,-14405.,-16226.
1420.000000000,-4707.0,-4436.0,-1682.3,-14405.,-16225.
1421.000000000,-4705.4,-4435.2,-1681.9,-14404.,-16225.
1422.000000000,-4703.8,-4434.4,-1681.5,-14404.,-16225.
1423.000000000,-4702.2,-4433.7,-1681.2,-14404.,-16224.
1424.000000000,-4700.7,-4433.0,-1680.8,-14404.,-16224.
1425.000000000,-4699.1,-4432.3,-1680.5,-14404.,-16224.
1426.000000000,-4698.1,-4432.1,-1680.5,-14403.,-16224.
1427.000000000,-4696.7,-4431.4,-1680.2,-14403.,-16223.
1428.000000000,-4695.3,-4430.6,-1679.8,-14403.,-16223.
1429.000000000,-4693.8,-4429.9,-1679.5,-14403.,-16223.
1430.000000000,-4692.3,-4429.2,-1679.1,-14403.,-16223.
1431.000000000,-4690.8,-4428.5,-1678.8,-14402.,-16222.
1432.000000000,-4689.3,-4427.8,-1678.5,-14402.,-16222.
1433.000000000,-4689.9,-4429.5,-1679.8,-14402.,-16222.
1434.000000000,-4692.5,-4432.8,-1682.2,-14402.,-16221.
1435.000000000,-4703.9,-4445.3,-1690.8,-14402.,-16221.
1436.000000000,-4707.3,-4444.0,-1690.7,-14401.,-16221.
1437.000000000,-4706.9,-4440.7,-1688.9,-14401.,-16221.
1438.000000000,-4705.3,-4438.0,-1687.3,-14401.,-16220.
1439.000000000,-4703.4,-4435.8,-1685.8,-14401.,-16220.
1440.000000000,-4701.4,-4434.1,-1684.6,-14401.,-16220.
1441.000000000,-4699.5,-4432.6,-1683.5,-14401.,-16219.
1442.000000000,-4697.6,-4431.3,-1682.6,-14400.,-16219.
1443.000000000,-4696.0,-4430.4,-1682.0,-14400.,-16219.
1444.000000000,-4694.3,-4429.3,-1681.3,-14400.,-16219.
1445.000000000,-4692.6,-4428.2,-1680.6,-14400.,-16218.
1446.000000000,-4690.9,-4427.3,-1680.0,-14400.,-16218.
1447.000000000,-4689.2,-4426.4,-1679.5,-14399.,-16218.
1448.000000000,-4687.6,-4425.5,-1678.9,-14399.,-16218.
1449.000000000,-4685.9,-4424.7,-1678.4,-14399.,-16217.
1450.000000000,-4684.3,-4423.8,-1678.0,-14399.,-16217.
1451.000000000,-4682.7,-4423.0,-1677.5,-14399.,-16217.
1452.000000000,-4681.4,-4422.6,-1677.3,-14398.,-16216.
1453.000000000,-4679.9,-4421.8,-1676.9,-14398.,-16216.
1454.000000000,-4678.9,-4421.6,-1676.9,-14398.,-16216.
1455.000000000,-4677.5,-4420.8,-1676.5,-14398.,-16216.
1456.000000000,-4676.0,-4420.0,-1676.1,-14398.,-16215.
1457.000000000,-4674.4,-4419.2,-1675.7,-14397.,-16215.
1458.000000000,-4672.9,-4418.5,-1675.3,-14397.,-16215.
1459.000000000,-4671.4,-4417.7,-1675.0,-14397.,-16214.
1460.000000000,-4670.0,-4417.2,-1674.7,-14397.,-16214.
1461.000000000,-4668.6,-4416.5,-1674.4,-14397.,-16214.
1462.000000000,-4667.1,-4415.8,-1674.0,-14397.,-16214.
1463.000000000,-4665.9,-4415.4,-1673.9,-14396.,-16213.
1464.000000000,-4664.6,-4414.7,-1673.6,-14396.,-16213.
1465.000000000,-4663.1,-4414.0,-1673.3,-14396.,-16213.
1466.000000000,-4661.7,-4413.3,-1673.0,-14396.,-16213.
1467.000000000,-4660.3,-4412.6,-1672.6,-14396.,-16212.
1468.000000000,-4658.8,-4411.9,-1672.3,-14395.,-16212.
1469.000000000,-4657.4,-4411.3,-1672.0,-14395.,-16212.
1470.000000000,-4656.0,-4410.6,-1671.7,-14395.,-16211.
1471.000000000,-4654.6,-4410.0,-1671.5,-14395.,-16211.
1472.000000000,-4653.2,-4409.3,-1671.2,-14395.,-16211.
1473.000000000,-4651.8,-4408.7,-1670.9,-14394.,-16211.
1474.000000000,-4650.4,-4408.1,-1670.6,-14394.,-16210.
1475.000000000,-4649.5,-4408.0,-1670.7,-14394.,-16210.
1476.000000000,-4649.1,-4408.3,-1671.1,-14394.,-16210.
1477.000000000,-4650.0,-4409.8,-1672.3,-14394.,-16209.
1478.000000000,-4649.2,-4408.8,-1671.9,-14393.,-16209.
1479.000000000,-4650.4,-4410.7,-1673.3,-14393.,-16209.
1480.000000000,-4649.8,-4409.4,-1672.8,-14393.,-16209.
1481.000000000,-4648.5,-4408.2,-1672.1,-14393.,-16208.
1482.000000000,-4647.1,-4407.1,-1671.5,-14393.,-16208.
1483.000000000,-4645.6,-4406.1,-1670.9,-14392.,-16208.
1484.000000000,-4644.1,-4405.2,-1670.4,-14392.,-16208.
1485.000000000,-4642.7,-4404.4,-1670.0,-14392.,-16207.
1486.000000000,-4641.2,-4403.6,-1669.6,-14392.,-16207.
1487.000000000,-4639.8,-4402.9,-1669.2,-14392.,-16207.
1488.000000000,-4638.4,-4402.2,-1668.8,-14392.,-16206.
1489.000000000,-4637.1,-4401.6,-1668.6,-14391.,-16206.
1490.000000000,-4635.8,-4400.9,-1668.3,-14391.,-16206.
1491.000000000,-4634.4,-4400.3,-1667.9,-14391.,-16206.
1492.000000000,-4633.1,-4399.6,-1667.6,-14391.,-16205.
1493.000000000,-4631.7,-4398.9,-1667.3,-14391.,-16205.
1494.000000000,-4630.4,-4398.3,-1667.0,-14390.,-16205.
1495.000000000,-4629.1,-4397.6,-1666.7,-14390.,-16205.
1496.000000000,-4627.7,-4397.0,-1666.4,-14390.,-16204.
1497.000000000,-4626.5,-4396.5,-1666.2,-14390.,-16204.
1498.000000000,-4625.2,-4395.8,-1666.0,-14390.,-16204.
1499.000000000,-4623.9,-4395.2,-1665.7,-14389.,-16203.
1500.000000000,-4622.6,-4394.6,-1665.4,-14389.,-16203.
1501.000000000,-4621.3,-4394.0,-1665.2,-14389.,-16203.
1502.000000000,-4620.1,-4393.3,-1664.9,-14389.,-16203.
1503.000000000,-4618.8,-4392.7,-1664.6,-14389.,-16202.
1504.000000000,-4617.5,-4392.1,-1664.4,-14388.,-16202.
1505.000000000,-4616.2,-4391.5,-1664.2,-14388.,-16202.
1506.000000000,-4622.8,-4400.4,-1670.1,-14388.,-16201.
1507.000000000,-4624.0,-4399.0,-1669.7,-14388.,-16201.
1508.000000000,-4623.3,-4397.0,-1668.8,-14388.,-16201.
1509.000000000,-4622.1,-4395.7,-1668.0,-14388.,-16201.
1510.000000000,-4620.7,-4394.4,-1667.2,-14387.,-16200.
1511.000000000,-4619.2,-4393.2,-1666.5,-14387.,-16200.
1512.000000000,-4618.8,-4393.5,-1666.8,-14387.,-16200.
1513.000000000,-4617.6,-4392.5,-1666.2,-14387.,-16200.
1514.000000000,-4616.3,-4391.5,-1665.6,-14387.,-16199.
1515.000000000,-4614.9,-4390.5,-1665.1,-14386.,-16199.
1516.000000000,-4613.4,-4389.7,-1664.6,-14386.,-16199.
1517.000000000,-4612.1,-4388.9,-1664.2,-14386.,-16198.
1518.000000000,-4610.7,-4388.1,-1663.8,-14386.,-16198.
1519.000000000,-4609.3,-4387.4,-1663.4,-14386.,-16198.
1520.000000000,-4608.0,-4386.7,-1663.0,-14385.,-16198.
1521.000000000,-4606.6,-4386.0,-1662.7,-14385.,-16197.
1522.000000000,-4605.3,-4385.4,-1662.3,-14385.,-16197.
1523.000000000,-4604.0,-4384.7,-1662.0,-14385.,-16197.
1524.000000000,-4602.7,-4384.1,-1661.7,-14385.,-16197.
1525.000000000,-4602.0,-4384.1,-1661.9,-14384.,-16196.
1526.000000000,-4600.8,-4383.4,-1661.6,-14384.,-16196.
1527.000000000,-4599.6,-4382.7,-1661.2,-14384.,-16196.
1528.000000000,-4598.3,-4382.0,-1660.9,-14384.,-16195.
1529.000000000,-4597.1,-4381.4,-1660.6,-14384.,-16195.
1530.000000000,-4595.8,-4380.7,-1660.3,-14383.,-16195.
1531.000000000,-4594.7,-4380.3,-1660.1,-14383.,-16195.
1532.000000000,-4593.5,-4379.6,-1659.9,-14383.,-16194.
1533.000000000,-4592.2,-4379.0,-1659.6,-14383.,-16194.
1534.000000000,-4591.0,-4378.4,-1659.3,-14383.,-16194.
1535.000000000,-4589.8,-4377.8,-1659.1,-14383.,-16194.
1536.000000000,-4588.5,-4377.2,-1658.8,-14382.,-16193.
1537.000000000,-4587.3,-4376.6,-1658.5,-14382.,-16193.
1538.000000000,-4586.1,-4376.0,-1658.3,-14382.,-16193.
1539.000000000,-4584.9,-4375.4,-1658.1,-14382.,-16193.
1540.000000000,-4583.7,-4374.8,-1657.8,-14382.,-16192.
1541.000000000,-4582.5,-4374.3,-1657.6,-14381.,-16192.
1542.000000000,-4581.3,-4373.7,-1657.3,-14381.,-16192.
1543.000000000,-4580.1,-4373.1,-1657.1,-14381.,-16191.
1544.000000000,-4579.0,-4372.7,-1656.9,-14381.,-16191.
1545.000000000,-4577.8,-4372.1,-1656.7,-14381.,-16191.
1546.000000000,-4576.7,-4371.5,-1656.5,-14380.,-16191.
1547.000000000,-4575.5,-4370.9,-1656.2,-14380.,-16190.
1548.000000000,-4574.3,-4370.4,-1656.0,-14380.,-16190.
1549.000000000,-4576.6,-4374.0,-1658.5,-14380.,-16190.
1550.000000000,-4576.5,-4373.0,-1658.2,-14380.,-16190.
1551.000000000,-4575.6,-4371.9,-1657.7,-14379.,-16189.
1552.000000000,-4574.4,-4370.9,-1657.2,-14379.,-16189.
1553.000000000,-4579.8,-4378.0,-1661.9,-14379.,-16189.
1554.000000000,-4580.5,-4376.5,-1661.4,-14379.,-16188.
1555.000000000,-4579.7,-4374.7,-1660.5,-14379.,-16188.
1556.000000000,-4578.4,-4373.2,-1659.6,-14379.,-16188.
1557.000000000,-4577.0,-4371.9,-1658.8,-14378.,-16188.
1558.000000000,-4575.6,-4370.9,-1658.1,-14378.,-16187.
1559.000000000,-4574.2,-4369.9,-1657.5,-14378.,-16187.
1560.000000000,-4572.8,-4369.0,-1657.0,-14378.,-16187.
1561.000000000,-4571.5,-4368.2,-1656.5,-14378.,-16187.
1562.000000000,-4572.3,-4370.0,-1657.8,-14377.,-16186.
1563.000000000,-4572.2,-4369.8,-1657.8,-14377.,-16186.
1564.000000000,-4572.0,-4369.5,-1657.8,-14377.,-16186.
1565.000000000,-4573.9,-4371.9,-1659.5,-14377.,-16185.
1566.000000000,-4573.5,-4370.6,-1658.8,-14377.,-16185.
1567.000000000,-4572.6,-4369.4,-1658.2,-14376.,-16185.
1568.000000000,-4572.3,-4369.4,-1658.3,-14376.,-16185.
1569.000000000,-4571.2,-4368.2,-1657.6,-14376.,-16184.
1570.000000000,-4569.8,-4367.1,-1656.9,-14376.,-16184.
1571.000000000,-4568.4,-4366.1,-1656.3,-14376.,-16184.
1572.000000000,-4567.0,-4365.2,-1655.7,-14376.,-16184.
1573.000000000,-4565.7,-4364.4,-1655.2,-14375.,-16183.
1574.000000000,-4564.3,-4363.6,-1654.8,-14375.,-16183.
1575.000000000,-4563.0,-4362.9,-1654.4,-14375.,-16183.
1576.000000000,-4561.6,-4362.1,-1654.0,-14375.,-16182.
1577.000000000,-4560.3,-4361.5,-1653.6,-14375.,-16182.
1578.000000000,-4559.1,-4360.8,-1653.3,-14374.,-16182.
1579.000000000,-4557.8,-4360.1,-1652.9,-14374.,-16182.
1580.000000000,-4556.5,-4359.5,-1652.6,-14374.,-16181.
1581.000000000,-4555.3,-4358.9,-1652.3,-14374.,-16181.
1582.000000000,-4554.0,-4358.3,-1652.0,-14374.,-16181.
1583.000000000,-4552.8,-4357.7,-1651.7,-14373.,-16181.
1584.000000000,-4551.5,-4357.1,-1651.4,-14373.,-16180.
1585.000000000,-4550.3,-4356.5,-1651.2,-14373.,-16180.
1586.000000000,-4549.1,-4355.9,-1650.9,-14373.,-16180.
1587.000000000,-4547.9,-4355.3,-1650.6,-14373.,-16180.
1588.000000000,-4546.7,-4354.7,-1650.4,-14372.,-16179.
1589.000000000,-4545.5,-4354.2,-1650.1,-14372.,-16179.
1590.000000000,-4544.3,-4353.6,-1649.9,-14372.,-16179.
1591.000000000,-4543.1,-4353.1,-1649.6,-14372.,-16178.
1592.000000000,-4544.7,-4355.8,-1651.6,-14372.,-16178.
1593.000000000,-4544.3,-4354.9,-1651.3,-14372.,-16178.
1594.000000000,-4543.4,-4353.9,-1650.8,-14371.,-16178.
1595.000000000,-4542.2,-4353.0,-1650.3,-14371.,-16177.
1596.000000000,-4541.0,-4352.2,-1649.9,-14371.,-16177.
1597.000000000,-4539.7,-4351.5,-1649.5,-14371.,-16177.
1598.000000000,-4538.6,-4350.9,-1649.3,-14371.,-16177.
1599.000000000,-4537.4,-4350.3,-1648.9,-14370.,-16176.
1600.000000000,-4536.2,-4349.6,-1648.6,-14370.,-16176.
1601.000000000,-4540.3,-4355.4,-1652.5,-14370.,-16176.
1602.000000000,-4541.1,-4354.7,-1652.5,-14370.,-16176.
1603.000000000,-4544.8,-4358.5,-1655.2,-14370.,-16175.
1604.000000000,-4545.0,-4356.8,-1654.4,-14369.,-16175.
1605.000000000,-4544.2,-4355.1,-1653.5,-14369.,-16175.
1606.000000000,-4542.9,-4353.6,-1652.5,-14369.,-16174.
1607.000000000,-4541.4,-4352.3,-1651.7,-14369.,-16174.
1608.000000000,-4540.0,-4351.2,-1651.0,-14369.,-16174.
1609.000000000,-4538.5,-4350.3,-1650.4,-14369.,-16174.
1610.000000000,-4542.5,-4355.8,-1654.0,-14368.,-16173.
1611.000000000,-4542.9,-4354.6,-1653.5,-14368.,-16173.
1612.000000000,-4559.5,-4374.0,-1666.4,-14368.,-16173.
1613.000000000,-4565.5,-4373.2,-1666.9,-14368.,-16173.
1614.000000000,-4566.3,-4369.4,-1664.8,-14368.,-16172.
1615.000000000,-4566.2,-4367.2,-1663.4,-14367.,-16172.
1616.000000000,-4567.7,-4367.9,-1663.8,-14367.,-16172.
1617.000000000,-4567.0,-4365.6,-1662.3,-14367.,-16172.
1618.000000000,-4565.3,-4363.1,-1660.5,-14367.,-16171.
1619.000000000,-4563.4,-4361.0,-1658.8,-14367.,-16171.
1620.000000000,-4561.4,-4359.2,-1657.5,-14366.,-16171.
1621.000000000,-4559.4,-4357.7,-1656.3,-14366.,-16170.
1622.000000000,-4557.6,-4356.3,-1655.2,-14366.,-16170.
1623.000000000,-4555.8,-4355.1,-1654.3,-14366.,-16170.
1624.000000000,-4554.0,-4354.0,-1653.5,-14366.,-16170.
1625.000000000,-4552.3,-4353.0,-1652.7,-14366.,-16169.
1626.000000000,-4550.6,-4352.0,-1652.0,-14365.,-16169.
1627.000000000,-4549.0,-4351.1,-1651.4,-14365.,-16169.
1628.000000000,-4547.4,-4350.3,-1650.9,-14365.,-16169.
1629.000000000,-4545.9,-4349.5,-1650.3,-14365.,-16168.
1630.000000000,-4544.3,-4348.7,-1649.8,-14365.,-16168.
1631.000000000,-4542.8,-4347.9,-1649.4,-14364.,-16168.
1632.000000000,-4541.3,-4347.2,-1648.9,-14364.,-16168.
1633.000000000,-4539.8,-4346.5,-1648.5,-14364.,-16167.
1634.000000000,-4538.3,-4345.8,-1648.1,-14364.,-16167.
1635.000000000,-4536.8,-4345.1,-1647.7,-14364.,-16167.
1636.000000000,-4535.5,-4344.5,-1647.4,-14363.,-16167.
1637.000000000,-4534.0,-4343.8,-1647.0,-14363.,-16166.
1638.000000000,-4532.7,-4343.2,-1646.7,-14363.,-16166.
1639.000000000,-4532.7,-4344.4,-1647.5,-14363.,-16166.
1640.000000000,-4532.1,-4343.9,-1647.4,-14363.,-16165.
1641.000000000,-4530.9,-4343.0,-1647.0,-14363.,-16165.
1642.000000000,-4529.5,-4342.2,-1646.5,-14362.,-16165.
1643.000000000,-4528.1,-4341.4,-1646.1,-14362.,-16165.
1644.000000000,-4526.7,-4340.7,-1645.7,-14362.,-16164.
1645.000000000,-4525.3,-4340.0,-1645.3,-14362.,-16164.
1646.000000000,-4523.9,-4339.4,-1645.0,-14362.,-16164.
1647.000000000,-4522.7,-4338.9,-1644.8,-14361.,-16164.
1648.000000000,-4521.6,-4338.5,-1644.6,-14361.,-16163.
1649.000000000,-4522.4,-4340.3,-1645.9,-14361.,-16163.
1650.000000000,-4524.3,-4342.6,-1647.6,-14361.,-16163.
1651.000000000,-4523.9,-4341.3,-1647.0,-14361.,-16163.
1652.000000000,-4522.7,-4340.0,-1646.3,-14360.,-16162.
1653.000000000,-4521.3,-4338.9,-1645.7,-14360.,-16162.
1654.000000000,-4519.9,-4337.9,-1645.1,-14360.,-16162.
1655.000000000,-4518.5,-4337.1,-1644.6,-14360.,-16161.
1656.000000000,-4517.5,-4336.8,-1644.5,-14360.,-16161.
1657.000000000,-4517.1,-4337.2,-1644.8,-14360.,-16161.
1658.000000000,-4517.5,-4338.1,-1645.5,-14359.,-16161.
1659.000000000,-4517.3,-4337.8,-1645.5,-14359.,-16160.
1660.000000000,-4516.6,-4337.1,-1645.2,-14359.,-16160.
1661.000000000,-4515.6,-4336.3,-1644.8,-14359.,-16160.
1662.000000000,-4514.3,-4335.3,-1644.2,-14359.,-16160.
1663.000000000,-4512.9,-4334.4,-1643.6,-14358.,-16159.
1664.000000000,-4511.5,-4333.6,-1643.2,-14358.,-16159.
1665.000000000,-4510.1,-4332.8,-1642.7,-14358.,-16159.
1666.000000000,-4513.8,-4338.3,-1646.4,-14358.,-16159.
1667.000000000,-4514.1,-4337.1,-1645.9,-14358.,-16158.
1668.000000000,-4513.1,-4335.6,-1645.1,-14358.,-16158.
1669.000000000,-4511.7,-4334.3,-1644.3,-14357.,-16158.
1670.000000000,-4510.3,-4333.2,-1643.7,-14357.,-16158.
1671.000000000,-4508.8,-4332.2,-1643.1,-14357.,-16157.
1672.000000000,-4507.3,-4331.4,-1642.5,-14357.,-16157.
1673.000000000,-4506.5,-4331.3,-1642.5,-14357.,-16157.
1674.000000000,-4505.6,-4330.9,-1642.3,-14356.,-16157.
1675.000000000,-4505.2,-4331.1,-1642.6,-14356.,-16156.
1676.000000000,-4505.2,-4331.4,-1642.9,-14356.,-16156.
1677.000000000,-4504.2,-4330.4,-1642.4,-14356.,-16156.
1678.000000000,-4503.0,-4329.5,-1641.9,-14356.,-16155.
1679.000000000,-4501.6,-4328.6,-1641.4,-14355.,-16155.
1680.000000000,-4500.2,-4327.8,-1640.9,-14355.,-16155.
1681.000000000,-4499.2,-4327.4,-1640.7,-14355.,-16155.
1682.000000000,-4504.5,-4334.6,-1645.5,-14355.,-16154.
1683.000000000,-4505.2,-4333.2,-1645.0,-14355.,-16154.
1684.000000000,-4504.4,-4331.5,-1644.1,-14355.,-16154.
1685.000000000,-4503.0,-4330.0,-1643.2,-14354.,-16154.
1686.000000000,-4501.5,-4328.8,-1642.4,-14354.,-16153.
1687.000000000,-4500.0,-4327.7,-1641.7,-14354.,-16153.
1688.000000000,-4498.5,-4326.8,-1641.1,-14354.,-16153.
1689.000000000,-4497.6,-4326.5,-1640.9,-14354.,-16153.
1690.000000000,-4496.5,-4325.9,-1640.6,-14353.,-16152.
1691.000000000,-4495.2,-4325.0,-1640.1,-14353.,-16152.
1692.000000000,-4493.8,-4324.3,-1639.6,-14353.,-16152.
1693.000000000,-4492.5,-4323.5,-1639.2,-14353.,-16152.
1694.000000000,-4491.1,-4322.8,-1638.8,-14353.,-16151.
1695.000000000,-4489.8,-4322.1,-1638.4,-14352.,-16151.
1696.000000000,-4488.4,-4321.4,-1638.1,-14352.,-16151.
1697.000000000,-4488.7,-4322.7,-1639.0,-14352.,-16151.
1698.000000000,-4489.9,-4324.3,-1640.2,-14352.,-16150.
1699.000000000,-4489.6,-4323.5,-1639.9,-14352.,-16150.
1700.000000000,-4489.7,-4323.9,-1640.3,-14352.,-16150.
1701.000000000,-4488.8,-4322.8,-1639.7,-14351.,-16150.
1702.000000000,-4487.5,-4321.7,-1639.1,-14351.,-16149.
1703.000000000,-4486.1,-4320.7,-1638.5,-14351.,-16149.
1704.000000000,-4484.7,-4319.8,-1638.0,-14351.,-16149.
1705.000000000,-4483.4,-4319.1,-1637.5,-14351.,-16148.
1706.000000000,-4482.0,-4318.3,-1637.1,-14350.,-16148.
1707.000000000,-4480.7,-4317.6,-1636.7,-14350.,-16148.
1708.000000000,-4479.4,-4317.1,-1636.4,-14350.,-16148.
1709.000000000,-4478.2,-4316.4,-1636.0,-14350.,-16147.
1710.000000000,-4476.9,-4315.8,-1635.7,-14350.,-16147.
1711.000000000,-4475.7,-4315.2,-1635.4,-14350.,-16147.
1712.000000000,-4474.4,-4314.6,-1635.1,-14349.,-16147.
1713.000000000,-4473.1,-4314.0,-1634.8,-14349.,-16146.
1714.000000000,-4471.9,-4313.4,-1634.5,-14349.,-16146.
1715.000000000,-4470.7,-4312.8,-1634.3,-14349.,-16146.
1716.000000000,-4469.5,-4312.3,-1634.0,-14349.,-16146.
1717.000000000,-4468.2,-4311.7,-1633.7,-14348.,-16145.
1718.000000000,-4467.0,-4311.2,-1633.5,-14348.,-16145.
1719.000000000,-4465.8,-4310.6,-1633.3,-14348.,-16145.
1720.000000000,-4464.6,-4310.1,-1633.0,-14348.,-16145.
1721.000000000,-4463.5,-4309.5,-1632.8,-14348.,-16144.
1722.000000000,-4462.3,-4309.0,-1632.5,-14347.,-16144.
1723.000000000,-4461.1,-4308.5,-1632.3,-14347.,-16144.
1724.000000000,-4460.1,-4308.1,-1632.2,-14347.,-16144.
1725.000000000,-4459.0,-4307.6,-1632.0,-14347.,-16143.
1726.000000000,-4457.8,-4307.0,-1631.7,-14347.,-16143.
1727.000000000,-4456.8,-4306.6,-1631.6,-14347.,-16143.
1728.000000000,-4455.7,-4306.1,-1631.4,-14346.,-16143.
1729.000000000,-4460.2,-4312.4,-1635.7,-14346.,-16142.
1730.000000000,-4464.2,-4315.4,-1638.0,-14346.,-16142.
1731.000000000,-4476.0,-4327.4,-1646.4,-14346.,-16142.
1732.000000000,-4489.9,-4338.1,-1654.2,-14346.,-16142.
1733.000000000,-4498.0,-4339.7,-1656.1,-14345.,-16141.
1734.000000000,-4500.4,-4336.6,-1654.6,-14345.,-16141.
1735.000000000,-4500.0,-4332.8,-1652.1,-14345.,-16141.
1736.000000000,-4498.2,-4329.1,-1649.5,-14345.,-16141.
1737.000000000,-4496.0,-4326.2,-1647.3,-14345.,-16140.
1738.000000000,-4497.1,-4327.9,-1648.1,-14345.,-16140.
1739.000000000,-4496.6,-4326.3,-1646.9,-14344.,-16140.
1740.000000000,-4495.0,-4324.0,-1645.2,-14344.,-16139.
1741.000000000,-4493.0,-4322.1,-1643.7,-14344.,-16139.
1742.000000000,-4491.1,-4320.4,-1642.4,-14344.,-16139.
1743.000000000,-4489.2,-4318.9,-1641.3,-14344.,-16139.
1744.000000000,-4489.1,-4319.8,-1641.7,-14343.,-16138.
1745.000000000,-4487.9,-4318.5,-1640.8,-14343.,-16138.
1746.000000000,-4486.3,-4317.2,-1639.9,-14343.,-16138.
1747.000000000,-4484.6,-4315.9,-1639.0,-14343.,-16138.
1748.000000000,-4482.9,-4314.9,-1638.2,-14343.,-16137.
1749.000000000,-4481.2,-4313.9,-1637.5,-14343.,-16137.
1750.000000000,-4479.5,-4313.0,-1636.8,-14342.,-16137.
1751.000000000,-4477.9,-4312.1,-1636.3,-14342.,-16137.
1752.000000000,-4476.3,-4311.3,-1635.7,-14342.,-16136.
1753.000000000,-4474.8,-4310.5,-1635.2,-14342.,-16136.
1754.000000000,-4473.2,-4309.7,-1634.7,-14342.,-16136.
1755.000000000,-4471.7,-4309.0,-1634.2,-14341.,-16136.
1756.000000000,-4470.2,-4308.3,-1633.8,-14341.,-16135.
1757.000000000,-4468.7,-4307.6,-1633.4,-14341.,-16135.
1758.000000000,-4467.2,-4307.0,-1633.0,-14341.,-16135.
1759.000000000,-4465.7,-4306.3,-1632.7,-14341.,-16135.
1760.000000000,-4464.3,-4305.7,-1632.3,-14341.,-16134.
1761.000000000,-4462.9,-4305.1,-1632.0,-14340.,-16134.
1762.000000000,-4461.5,-4304.4,-1631.6,-14340.,-16134.
1763.000000000,-4460.1,-4303.8,-1631.3,-14340.,-16134.
1764.000000000,-4458.7,-4303.2,-1631.0,-14340.,-16133.
1765.000000000,-4457.3,-4302.7,-1630.7,-14340.,-16133.
1766.000000000,-4456.0,-4302.1,-1630.4,-14339.,-16133.
1767.000000000,-4454.6,-4301.5,-1630.2,-14339.,-16133.
1768.000000000,-4453.3,-4301.0,-1629.9,-14339.,-16132.
1769.000000000,-4451.9,-4300.4,-1629.6,-14339.,-16132.
1770.000000000,-4450.6,-4299.8,-1629.3,-14339.,-16132.
1771.000000000,-4449.3,-4299.3,-1629.1,-14338.,-16132.
1772.000000000,-4448.0,-4298.7,-1628.8,-14338.,-16131.
1773.000000000,-4446.7,-4298.2,-1628.6,-14338.,-16131.
1774.000000000,-4445.5,-4297.7,-1628.4,-14338.,-16131.
1775.000000000,-4444.2,-4297.2,-1628.1,-14338.,-16130.
1776.000000000,-4443.0,-4296.6,-1627.9,-14338.,-16130.
1777.000000000,-4442.2,-4296.7,-1628.1,-14337.,-16130.
1778.000000000,-4441.2,-4296.1,-1627.8,-14337.,-16130.
1779.000000000,-4440.1,-4295.7,-1627.6,-14337.,-16129.
1780.000000000,-4438.9,-4295.1,-1627.4,-14337.,-16129.
1781.000000000,-4437.7,-4294.5,-1627.1,-14337.,-16129.
1782.000000000,-4436.4,-4293.9,-1626.8,-14337.,-16128.
1783.000000000,-4435.2,-4293.3,-1626.6,-14336.,-16128.
1784.000000000,-4434.0,-4292.8,-1626.3,-14336.,-16128.
1785.000000000,-4432.8,-4292.3,-1626.1,-14336.,-16127.
1786.000000000,-4431.6,-4291.7,-1625.9,-14336.,-16127.
1787.000000000,-4430.4,-4291.2,-1625.6,-14336.,-16127.
1788.000000000,-4429.2,-4290.7,-1625.4,-14335.,-16127.
1789.000000000,-4428.0,-4290.2,-1625.2,-14335.,-16126.
1790.000000000,-4426.8,-4289.6,-1625.0,-14335.,-16126.
1791.000000000,-4425.7,-4289.1,-1624.8,-14335.,-16126.
1792.000000000,-4424.5,-4288.6,-1624.6,-14335.,-16125.
1793.000000000,-4423.4,-4288.1,-1624.4,-14335.,-16125.
1794.000000000,-4422.2,-4287.6,-1624.2,-14334.,-16125.
1795.000000000,-4421.1,-4287.1,-1624.0,-14334.,-16125.
1796.000000000,-4419.9,-4286.6,-1623.8,-14334.,-16124.
1797.000000000,-4418.8,-4286.1,-1623.6,-14334.,-16124.
1798.000000000,-4417.7,-4285.6,-1623.4,-14334.,-16124.
1799.000000000,-4416.6,-4285.1,-1623.2,-14334.,-16123.
1800.000000000,-4415.5,-4284.6,-1623.0,-14333.,-16123.
1801.000000000,-4415.9,-4286.0,-1624.0,-14333.,-16123.
1802.000000000,-4420.9,-4292.1,-1628.2,-14333.,-16123.
1803.000000000,-4423.1,-4292.6,-1629.1,-14333.,-16122.
1804.000000000,-4422.9,-4290.9,-1628.2,-14333.,-16122.
1805.000000000,-4421.8,-4289.3,-1627.3,-14332.,-16122.
1806.000000000,-4420.5,-4288.0,-1626.5,-14332.,-16122.
1807.000000000,-4419.2,-4286.9,-1625.8,-14332.,-16121.
1808.000000000,-4417.9,-4286.0,-1625.3,-14332.,-16121.
1809.000000000,-4416.6,-4285.2,-1624.7,-14332.,-16121.
1810.000000000,-4415.3,-4284.4,-1624.3,-14332.,-16120.
1811.000000000,-4414.3,-4284.0,-1624.0,-14331.,-16120.
1812.000000000,-4415.1,-4285.7,-1625.2,-14331.,-16120.
1813.000000000,-4414.5,-4284.8,-1624.8,-14331.,-16120.
1814.000000000,-4413.8,-4284.3,-1624.6,-14331.,-16119.
1815.000000000,-4412.8,-4283.4,-1624.1,-14331.,-16119.
1816.000000000,-4411.6,-4282.6,-1623.7,-14330.,-16119.
1817.000000000,-4410.3,-4281.8,-1623.2,-14330.,-16118.
1818.000000000,-4409.2,-4281.2,-1622.9,-14330.,-16118.
1819.000000000,-4408.0,-4280.5,-1622.5,-14330.,-16118.
1820.000000000,-4406.8,-4279.9,-1622.2,-14330.,-16118.
1821.000000000,-4405.6,-4279.2,-1621.8,-14330.,-16117.
1822.000000000,-4404.7,-4278.9,-1621.7,-14329.,-16117.
1823.000000000,-4403.7,-4278.5,-1621.5,-14329.,-16117.
1824.000000000,-4402.6,-4277.9,-1621.2,-14329.,-16116.
1825.000000000,-4401.5,-4277.3,-1621.0,-14329.,-16116.
1826.000000000,-4400.4,-4276.7,-1620.7,-14329.,-16116.
1827.000000000,-4399.3,-4276.2,-1620.4,-14329.,-16116.
1828.000000000,-4398.2,-4275.7,-1620.2,-14328.,-16115.
1829.000000000,-4397.1,-4275.1,-1620.0,-14328.,-16115.
1830.000000000,-4396.0,-4274.6,-1619.7,-14328.,-16115.
1831.000000000,-4394.9,-4274.1,-1619.5,-14328.,-16115.
1832.000000000,-4393.9,-4273.6,-1619.3,-14328.,-16114.
1833.000000000,-4392.8,-4273.1,-1619.0,-14327.,-16114.
1834.000000000,-4391.7,-4272.5,-1618.8,-14327.,-16114.
1835.000000000,-4390.6,-4272.0,-1618.6,-14327.,-16113.
1836.000000000,-4389.6,-4271.5,-1618.4,-14327.,-16113.
1837.000000000,-4388.5,-4271.1,-1618.2,-14327.,-16113.
1838.000000000,-4387.5,-4270.6,-1618.0,-14327.,-16113.
1839.000000000,-4386.4,-4270.1,-1617.8,-14326.,-16112.
1840.000000000,-4385.4,-4269.6,-1617.6,-14326.,-16112.
1841.000000000,-4384.4,-4269.1,-1617.4,-14326.,-16112.
1842.000000000,-4383.4,-4268.8,-1617.3,-14326.,-16111.
1843.000000000,-4382.5,-4268.3,-1617.1,-14326.,-16111.
1844.000000000,-4381.4,-4267.8,-1616.9,-14326.,-16111.
1845.000000000,-4380.5,-4267.4,-1616.8,-14325.,-16111.
1846.000000000,-4379.6,-4267.0,-1616.6,-14325.,-16110.
1847.000000000,-4378.6,-4266.5,-1616.4,-14325.,-16110.
1848.000000000,-4377.6,-4266.0,-1616.2,-14325.,-16110.
1849.000000000,-4376.6,-4265.5,-1616.0,-14325.,-16110.
1850.000000000,-4375.6,-4265.0,-1615.9,-14324.,-16109.
1851.000000000,-4374.6,-4264.5,-1615.7,-14324.,-16109.
1852.000000000,-4373.6,-4264.0,-1615.5,-14324.,-16109.
1853.000000000,-4372.6,-4263.6,-1615.3,-14324.,-16108.
1854.000000000,-4371.7,-4263.1,-1615.1,-14324.,-16108.
1855.000000000,-4370.7,-4262.6,-1614.9,-14324.,-16108.
1856.000000000,-4369.7,-4262.2,-1614.8,-14323.,-16108.
1857.000000000,-4368.8,-4261.7,-1614.6,-14323.,-16107.
1858.000000000,-4367.8,-4261.2,-1614.4,-14323.,-16107.
1859.000000000,-4366.8,-4260.8,-1614.2,-14323.,-16107.
1860.000000000,-4366.0,-4260.5,-1614.1,-14323.,-16107.
1861.000000000,-4365.1,-4260.0,-1614.0,-14323.,-16106.
1862.000000000,-4364.1,-4259.5,-1613.8,-14322.,-16106.
1863.000000000,-4363.2,-4259.0,-1613.6,-14322.,-16106.
1864.000000000,-4362.3,-4258.6,-1613.5,-14322.,-16106.
1865.000000000,-4361.4,-4258.2,-1613.3,-14322.,-16105.
1866.000000000,-4360.5,-4257.7,-1613.1,-14322.,-16105.
1867.000000000,-4359.5,-4257.2,-1612.9,-14321.,-16105.
1868.000000000,-4358.6,-4256.8,-1612.8,-14321.,-16104.
1869.000000000,-4357.7,-4256.3,-1612.6,-14321.,-16104.
1870.000000000,-4357.1,-4256.3,-1612.7,-14321.,-16104.
1871.000000000,-4356.4,-4256.0,-1612.6,-14321.,-16104.
1872.000000000,-4355.6,-4255.5,-1612.4,-14321.,-16103.
1873.000000000,-4354.7,-4254.9,-1612.2,-14320.,-16103.
1874.000000000,-4353.8,-4254.4,-1612.0,-14320.,-16103.
1875.000000000,-4352.8,-4254.0,-1611.8,-14320.,-16103.
1876.000000000,-4352.5,-4254.2,-1612.1,-14320.,-16102.
1877.000000000,-4353.3,-4255.6,-1613.2,-14320.,-16102.
1878.000000000,-4359.4,-4262.7,-1618.0,-14320.,-16102.
1879.000000000,-4361.0,-4261.8,-1618.0,-14319.,-16101.
1880.000000000,-4360.7,-4260.0,-1617.0,-14319.,-16101.
1881.000000000,-4359.8,-4258.6,-1616.2,-14319.,-16101.
1882.000000000,-4358.7,-4257.4,-1615.5,-14319.,-16101.
1883.000000000,-4357.6,-4256.3,-1614.8,-14319.,-16100.
1884.000000000,-4356.4,-4255.4,-1614.2,-14318.,-16100.
1885.000000000,-4355.3,-4254.6,-1613.7,-14318.,-16100.
1886.000000000,-4354.5,-4254.3,-1613.5,-14318.,-16100.
1887.000000000,-4353.5,-4253.6,-1613.1,-14318.,-16099.
1888.000000000,-4352.5,-4252.9,-1612.7,-14318.,-16099.
1889.000000000,-4351.4,-4252.2,-1612.3,-14318.,-16099.
1890.000000000,-4350.4,-4251.6,-1612.0,-14317.,-16099.
1891.000000000,-4349.3,-4251.0,-1611.7,-14317.,-16098.
1892.000000000,-4348.3,-4250.4,-1611.4,-14317.,-16098.
1893.000000000,-4347.3,-4249.9,-1611.1,-14317.,-16098.
1894.000000000,-4346.3,-4249.4,-1610.8,-14317.,-16098.
1895.000000000,-4345.3,-4248.8,-1610.6,-14317.,-16097.
1896.000000000,-4344.3,-4248.3,-1610.3,-14316.,-16097.
1897.000000000,-4343.3,-4247.8,-1610.1,-14316.,-16097.
1898.000000000,-4342.4,-4247.3,-1609.9,-14316.,-16096.
1899.000000000,-4341.4,-4246.8,-1609.7,-14316.,-16096.
1900.000000000,-4340.5,-4246.4,-1609.4,-14316.,-16096.
1901.000000000,-4339.5,-4245.9,-1609.2,-14315.,-16096.
1902.000000000,-4338.6,-4245.4,-1609.0,-14315.,-16095.
1903.000000000,-4337.6,-4244.9,-1608.8,-14315.,-16095.
1904.000000000,-4336.7,-4244.5,-1608.6,-14315.,-16095.
1905.000000000,-4335.8,-4244.0,-1608.5,-14315.,-16095.
1906.000000000,-4334.8,-4243.6,-1608.3,-14315.,-16094.
1907.000000000,-4333.9,-4243.1,-1608.1,-14314.,-16094.
1908.000000000,-4333.0,-4242.6,-1607.9,-14314.,-16094.
1909.000000000,-4332.1,-4242.2,-1607.7,-14314.,-16094.
1910.000000000,-4331.2,-4241.7,-1607.5,-14314.,-16093.
1911.000000000,-4330.3,-4241.3,-1607.4,-14314.,-16093.
1912.000000000,-4329.4,-4240.9,-1607.2,-14314.,-16093.
1913.000000000,-4328.8,-4240.8,-1607.3,-14313.,-16093.
1914.000000000,-4328.0,-4240.3,-1607.1,-14313.,-16092.
1915.000000000,-4327.1,-4239.8,-1606.9,-14313.,-16092.
1916.000000000,-4326.2,-4239.3,-1606.7,-14313.,-16092.
1917.000000000,-4325.3,-4238.9,-1606.5,-14313.,-16091.
1918.000000000,-4324.4,-4238.4,-1606.3,-14313.,-16091.
1919.000000000,-4323.6,-4238.0,-1606.1,-14312.,-16091.
1920.000000000,-4322.7,-4237.5,-1605.9,-14312.,-16091.
1921.000000000,-4321.8,-4237.1,-1605.8,-14312.,-16090.
1922.000000000,-4320.9,-4236.6,-1605.6,-14312.,-16090.
1923.000000000,-4320.0,-4236.2,-1605.4,-14312.,-16090.
1924.000000000,-4319.2,-4235.8,-1605.3,-14311.,-16090.
1925.000000000,-4318.3,-4235.3,-1605.1,-14311.,-16089.
1926.000000000,-4317.4,-4234.9,-1604.9,-14311.,-16089.
1927.000000000,-4316.6,-4234.5,-1604.8,-14311.,-16089.
1928.000000000,-4315.7,-4234.0,-1604.6,-14311.,-16089.
1929.000000000,-4314.9,-4233.6,-1604.4,-14311.,-16088.
1930.000000000,-4314.2,-4233.4,-1604.4,-14310.,-16088.
1931.000000000,-4313.4,-4232.9,-1604.3,-14310.,-16088.
1932.000000000,-4312.6,-4232.5,-1604.1,-14310.,-16088.
1933.000000000,-4311.7,-4232.0,-1603.9,-14310.,-16087.
1934.000000000,-4310.9,-4231.6,-1603.7,-14310.,-16087.
1935.000000000,-4310.0,-4231.2,-1603.6,-14310.,-16087.
1936.000000000,-4309.2,-4230.7,-1603.4,-14309.,-16087.
1937.000000000,-4308.4,-4230.3,-1603.3,-14309.,-16086.
1938.000000000,-4307.7,-4230.0,-1603.2,-14309.,-16086.
1939.000000000,-4306.9,-4229.6,-1603.0,-14309.,-16086.
1940.000000000,-4306.1,-4229.2,-1602.9,-14309.,-16086.
1941.000000000,-4305.2,-4228.7,-1602.7,-14308.,-16085.
1942.000000000,-4305.5,-4229.6,-1603.4,-14308.,-16085.
1943.000000000,-4305.0,-4229.0,-1603.2,-14308.,-16085.
1944.000000000,-4304.2,-4228.4,-1602.9,-14308.,-16084.
1945.000000000,-4303.4,-4227.9,-1602.7,-14308.,-16084.
1946.000000000,-4302.5,-4227.4,-1602.5,-14308.,-16084.
1947.000000000,-4301.7,-4226.9,-1602.2,-14307.,-16084.
1948.000000000,-4300.9,-4226.4,-1602.0,-14307.,-16083.
1949.000000000,-4300.3,-4226.3,-1602.1,-14307.,-16083.
1950.000000000,-4306.9,-4234.8,-1607.8,-14307.,-16083.
1951.000000000,-4309.5,-4235.0,-1608.4,-14307.,-16083.
1952.000000000,-4309.6,-4233.1,-1607.5,-14307.,-16082.
1953.000000000,-4308.8,-4231.5,-1606.6,-14306.,-16082.
1954.000000000,-4307.7,-4230.3,-1605.8,-14306.,-16082.
1955.000000000,-4306.7,-4229.2,-1605.1,-14306.,-16082.
1956.000000000,-4305.6,-4228.4,-1604.5,-14306.,-16081.
1957.000000000,-4304.5,-4227.6,-1604.0,-14306.,-16081.
1958.000000000,-4303.5,-4226.9,-1603.6,-14306.,-16081.
1959.000000000,-4302.5,-4226.2,-1603.2,-14305.,-16081.
1960.000000000,-4301.5,-4225.6,-1602.8,-14305.,-16080.
1961.000000000,-4300.5,-4225.0,-1602.5,-14305.,-16080.
1962.000000000,-4299.6,-4224.5,-1602.2,-14305.,-16080.
1963.000000000,-4298.7,-4223.9,-1601.9,-14305.,-16080.
1964.000000000,-4297.8,-4223.5,-1601.7,-14304.,-16079.
1965.000000000,-4296.9,-4223.0,-1601.4,-14304.,-16079.
1966.000000000,-4296.7,-4223.3,-1601.7,-14304.,-16079.
1967.000000000,-4303.0,-4231.3,-1607.1,-14304.,-16079.
1968.000000000,-4304.5,-4230.2,-1606.8,-14304.,-16078.
1969.000000000,-4304.1,-4228.4,-1605.9,-14304.,-16078.
1970.000000000,-4303.2,-4227.0,-1605.0,-14303.,-16078.
1971.000000000,-4302.1,-4225.8,-1604.3,-14303.,-16078.
1972.000000000,-4300.9,-4224.9,-1603.6,-14303.,-16077.
1973.000000000,-4299.8,-4224.0,-1603.1,-14303.,-16077.
1974.000000000,-4298.8,-4223.3,-1602.6,-14303.,-16077.
1975.000000000,-4297.7,-4222.6,-1602.2,-14303.,-16077.
1976.000000000,-4296.7,-4221.9,-1601.8,-14302.,-16076.
1977.000000000,-4295.7,-4221.3,-1601.4,-14302.,-16076.
1978.000000000,-4294.7,-4220.8,-1601.1,-14302.,-16076.
1979.000000000,-4293.7,-4220.2,-1600.8,-14302.,-16076.
1980.000000000,-4292.7,-4219.7,-1600.5,-14302.,-16075.
1981.000000000,-4292.1,-4219.6,-1600.5,-14301.,-16075.
1982.000000000,-4291.3,-4219.1,-1600.2,-14301.,-16075.
1983.000000000,-4290.4,-4218.5,-1600.0,-14301.,-16075.
1984.000000000,-4289.4,-4218.0,-1599.7,-14301.,-16074.
1985.000000000,-4288.5,-4217.5,-1599.4,-14301.,-16074.
1986.000000000,-4287.6,-4217.0,-1599.2,-14301.,-16074.
1987.000000000,-4286.7,-4216.5,-1599.0,-14300.,-16074.
1988.000000000,-4285.8,-4216.1,-1598.7,-14300.,-16073.
1989.000000000,-4284.9,-4215.6,-1598.5,-14300.,-16073.
1990.000000000,-4284.0,-4215.1,-1598.3,-14300.,-16073.
1991.000000000,-4283.1,-4214.7,-1598.1,-14300.,-16073.
1992.000000000,-4282.2,-4214.3,-1597.9,-14300.,-16072.
1993.000000000,-4281.3,-4213.8,-1597.7,-14299.,-16072.
1994.000000000,-4280.4,-4213.4,-1597.5,-14299.,-16072.
1995.000000000,-4279.6,-4213.0,-1597.4,-14299.,-16072.
1996.000000000,-4279.2,-4213.1,-1597.6,-14299.,-16071.
1997.000000000,-4278.5,-4212.7,-1597.4,-14299.,-16071.
1998.000000000,-4277.7,-4212.2,-1597.2,-14299.,-16071.
1999.000000000,-4276.9,-4211.8,-1597.0,-14298.,-16071.
2000.000000000,-4276.1,-4211.3,-1596.8,-14298.,-16070.
2001.000000000,-4275.2,-4210.8,-1596.6,-14298.,-16070.
2002.000000000,-4274.3,-4210.4,-1596.4,-14298.,-16070.
2003.000000000,-4273.5,-4210.0,-1596.2,-14298.,-16070.
2004.000000000,-4272.6,-4209.5,-1596.0,-14298.,-16069.
2005.000000000,-4271.8,-4209.1,-1595.9,-14297.,-16069.
2006.000000000,-4271.0,-4208.7,-1595.7,-14297.,-16069.
2007.000000000,-4270.5,-4208.7,-1595.8,-14297.,-16069.
2008.000000000,-4269.8,-4208.3,-1595.7,-14297.,-16068.
2009.000000000,-4269.0,-4207.8,-1595.5,-14297.,-16068.
2010.000000000,-4268.2,-4207.3,-1595.3,-14296.,-16068.
2011.000000000,-4267.3,-4206.9,-1595.1,-14296.,-16068.
2012.000000000,-4267.2,-4207.4,-1595.5,-14296.,-16067.
2013.000000000,-4267.9,-4208.4,-1596.3,-14296.,-16067.
2014.000000000,-4270.5,-4211.4,-1598.4,-14296.,-16067.
2015.000000000,-4273.9,-4214.2,-1600.6,-14296.,-16067.
2016.000000000,-4275.5,-4214.4,-1601.0,-14295.,-16066.
2017.000000000,-4277.5,-4215.5,-1601.9,-14295.,-16066.
2018.000000000,-4277.3,-4213.8,-1601.0,-14295.,-16066.
2019.000000000,-4276.4,-4212.3,-1600.1,-14295.,-16066.
2020.000000000,-4275.3,-4211.0,-1599.3,-14295.,-16065.
2021.000000000,-4274.2,-4210.0,-1598.6,-14295.,-16065.
2022.000000000,-4273.0,-4209.1,-1598.0,-14294.,-16065.
2023.000000000,-4272.0,-4208.3,-1597.4,-14294.,-16065.
2024.000000000,-4270.9,-4207.6,-1596.9,-14294.,-16064.
2025.000000000,-4269.9,-4206.9,-1596.5,-14294.,-16064.
2026.000000000,-4268.9,-4206.3,-1596.1,-14294.,-16064.
2027.000000000,-4267.9,-4205.7,-1595.8,-14294.,-16064.
2028.000000000,-4266.9,-4205.2,-1595.5,-14293.,-16063.
2029.000000000,-4265.9,-4204.7,-1595.2,-14293.,-16063.
2030.000000000,-4265.0,-4204.1,-1594.9,-14293.,-16063.
2031.000000000,-4264.1,-4203.6,-1594.6,-14293.,-16063.
2032.000000000,-4263.1,-4203.1,-1594.3,-14293.,-16062.
2033.000000000,-4262.2,-4202.7,-1594.1,-14292.,-16062.
2034.000000000,-4261.3,-4202.2,-1593.9,-14292.,-16062.
2035.000000000,-4260.4,-4201.7,-1593.6,-14292.,-16062.
2036.000000000,-4259.5,-4201.3,-1593.4,-14292.,-16061.
2037.000000000,-4258.6,-4200.9,-1593.2,-14292.,-16061.
2038.000000000,-4264.9,-4209.2,-1598.8,-14292.,-16061.
2039.000000000,-4266.5,-4208.3,-1598.7,-14291.,-16061.
2040.000000000,-4266.2,-4206.6,-1597.8,-14291.,-16060.
2041.000000000,-4265.3,-4205.2,-1597.0,-14291.,-16060.
2042.000000000,-4264.2,-4204.1,-1596.3,-14291.,-16060.
2043.000000000,-4263.1,-4203.2,-1595.7,-14291.,-16060.
2044.000000000,-4262.0,-4202.4,-1595.2,-14291.,-16059.
2045.000000000,-4261.0,-4201.7,-1594.7,-14290.,-16059.
2046.000000000,-4260.0,-4201.1,-1594.3,-14290.,-16059.
2047.000000000,-4258.9,-4200.5,-1593.9,-14290.,-16059.
2048.000000000,-4258.0,-4199.9,-1593.6,-14290.,-16058.
2049.000000000,-4259.8,-4202.7,-1595.5,-14290.,-16058.
2050.000000000,-4261.5,-4204.2,-1596.7,-14290.,-16058.
2051.000000000,-4263.9,-4206.1,-1598.1,-14289.,-16058.
2052.000000000,-4264.4,-4205.5,-1597.9,-14289.,-16057.
2053.000000000,-4263.8,-4204.0,-1597.1,-14289.,-16057.
2054.000000000,-4262.8,-4202.8,-1596.3,-14289.,-16057.
2055.000000000,-4261.6,-4201.7,-1595.6,-14289.,-16057.
2056.000000000,-4260.5,-4200.9,-1595.0,-14289.,-16057.
2057.000000000,-4259.4,-4200.1,-1594.5,-14288.,-16056.
2058.000000000,-4258.9,-4200.1,-1594.5,-14288.,-16056.
2059.000000000,-4259.2,-4200.8,-1595.0,-14288.,-16056.
2060.000000000,-4258.5,-4200.0,-1594.5,-14288.,-16056.
2061.000000000,-4257.6,-4199.1,-1594.0,-14288.,-16055.
2062.000000000,-4256.5,-4198.4,-1593.6,-14288.,-16055.
2063.000000000,-4255.5,-4197.7,-1593.1,-14287.,-16055.
2064.000000000,-4254.5,-4197.1,-1592.8,-14287.,-16055.
2065.000000000,-4253.5,-4196.5,-1592.4,-14287.,-16054.
2066.000000000,-4252.5,-4196.0,-1592.1,-14287.,-16054.
2067.000000000,-4251.5,-4195.4,-1591.8,-14287.,-16054.
2068.000000000,-4250.5,-4194.9,-1591.5,-14286.,-16054.
2069.000000000,-4249.5,-4194.4,-1591.3,-14286.,-16053.
