time,EAST,NORTH,WEST,PATH
1.000000000000,5666.3,2572.1,2781.2,25290.
2.000000000000,5666.1,2572.0,2781.2,25290.
3.000000000000,5665.8,2571.9,2780.9,25289.
4.000000000000,5665.4,2571.8,2779.2,25289.
5.000000000000,5664.9,2571.6,2777.7,25289.
6.000000000000,5664.4,2571.3,2776.5,25288.
7.000000000000,5663.7,2571.0,2775.3,25288.
8.000000000000,5663.0,2570.7,2774.0,25287.
9.000000000000,5662.2,2570.3,2766.2,25286.
10.00000000000,5661.3,2569.9,2756.8,25286.
11.00000000000,5660.3,2569.4,2755.3,25285.
12.00000000000,5659.3,2568.9,2755.1,25284.
13.00000000000,5658.3,2568.4,2755.0,25283.
14.00000000000,5657.1,2567.8,2754.8,25283.
15.00000000000,5656.0,2567.1,2754.2,25282.
16.00000000000,5654.7,2566.5,2753.3,25281.
17.00000000000,5653.5,2565.8,2752.2,25280.
18.00000000000,5652.1,2565.0,2750.8,25279.
19.00000000000,5650.8,2564.3,2749.3,25278.
20.00000000000,5649.4,2563.5,2747.7,25277.
21.00000000000,5648.0,2562.6,2745.9,25276.
22.00000000000,5646.5,2561.8,2744.1,25275.
23.00000000000,5645.0,2560.9,2742.2,25275.
24.00000000000,5643.5,2560.0,2740.2,25274.
25.00000000000,5642.0,2559.0,2738.2,25273.
26.00000000000,5640.4,2558.1,2736.3,25272.
27.00000000000,5638.8,2557.1,2734.3,25271.
28.00000000000,5637.2,2556.1,2732.3,25270.
29.00000000000,5635.6,2555.1,2730.4,25269.
30.00000000000,5634.0,2554.1,2728.5,25268.
31.00000000000,5632.4,2553.1,2726.6,25267.
32.00000000000,5630.7,2552.0,2724.7,25266.
33.00000000000,5629.1,2551.0,2722.9,25265.
34.00000000000,5627.5,2550.0,2721.2,25264.
35.00000000000,5625.8,2548.9,2719.4,25263.
36.00000000000,5624.2,2547.9,2717.7,25262.
37.00000000000,5622.6,2546.8,2716.1,25261.
38.00000000000,5621.0,2545.8,2714.5,25260.
39.00000000000,5619.4,2544.7,2712.9,25259.
40.00000000000,5617.8,2543.7,2711.4,25258.
41.00000000000,5616.2,2542.6,2709.8,25257.
42.00000000000,5614.7,2541.6,2708.4,25256.
43.00000000000,5613.1,2540.6,2707.0,25256.
44.00000000000,5611.6,2539.6,2705.6,25255.
45.00000000000,5610.1,2538.6,2704.3,25254.
46.00000000000,5608.7,2537.7,2703.0,25253.
47.00000000000,5607.3,2536.7,2701.8,25252.
48.00000000000,5605.8,2535.8,2700.5,25251.
49.00000000000,5604.5,2534.9,2699.4,25251.
50.00000000000,5603.1,2534.0,2698.2,25250.
51.00000000000,5601.8,2533.1,2697.1,25249.
52.00000000000,5600.5,2532.2,2695.6,25248.
53.00000000000,5599.2,2531.3,2694.6,25248.
54.00000000000,5598.0,2530.5,2693.6,25247.
55.00000000000,5596.7,2529.6,2692.6,25246.
56.00000000000,5595.5,2528.8,2691.4,25245.
57.00000000000,5594.3,2528.0,2690.5,25245.
58.00000000000,5593.2,2527.2,2689.6,25244.
59.00000000000,5592.1,2526.4,2688.8,25243.
60.00000000000,5591.0,2525.7,2688.0,25243.
61.00000000000,5589.9,2524.9,2687.3,25242.
62.00000000000,5588.9,2524.2,2686.5,25242.
63.00000000000,5587.9,2523.5,2685.8,25241.
64.00000000000,5586.9,2522.8,2685.1,25240.
65.00000000000,5586.0,2522.1,2684.4,25240.
66.00000000000,5585.1,2521.5,2683.7,25239.
67.00000000000,5584.2,2520.8,2683.0,25239.
68.00000000000,5583.3,2520.2,2682.4,25238.
69.00000000000,5582.4,2519.6,2680.7,25238.
70.00000000000,5581.6,2519.0,2680.0,25237.
71.00000000000,5580.8,2518.4,2679.5,25237.
72.00000000000,5579.9,2517.8,2679.1,25236.
73.00000000000,5579.2,2517.3,2678.6,25236.
74.00000000000,5578.4,2516.7,2678.2,25235.
75.00000000000,5577.6,2516.2,2677.8,25235.
76.00000000000,5576.9,2515.7,2677.3,25234.
77.00000000000,5576.2,2515.2,2676.9,25234.
78.00000000000,5575.5,2514.7,2676.4,25234.
79.00000000000,5574.8,2514.2,2675.9,25233.
80.00000000000,5574.1,2513.7,2675.4,25233.
81.00000000000,5573.5,2513.2,2674.9,25232.
82.00000000000,5572.8,2512.8,2673.8,25232.
83.00000000000,5572.2,2512.3,2673.3,25231.
84.00000000000,5571.6,2511.9,2672.9,25231.
85.00000000000,5571.0,2511.4,2672.6,25231.
86.00000000000,5570.4,2511.0,2672.2,25230.
87.00000000000,5569.8,2510.6,2671.9,25230.
88.00000000000,5569.2,2510.2,2671.5,25229.
89.00000000000,5568.7,2509.8,2671.2,25229.
90.00000000000,5568.1,2509.4,2670.8,25229.
91.00000000000,5567.6,2509.0,2670.5,25228.
92.00000000000,5567.1,2508.6,2670.1,25228.
93.00000000000,5566.6,2508.2,2667.0,25228.
94.00000000000,5566.1,2507.9,2666.5,25227.
95.00000000000,5565.6,2507.5,2666.4,25227.
96.00000000000,5565.1,2507.2,2666.5,25227.
97.00000000000,5564.6,2506.8,2666.6,25226.
98.00000000000,5564.2,2506.5,2666.6,25226.
99.00000000000,5563.7,2506.1,2666.5,25226.
100.0000000000,5563.3,2505.8,2666.4,25225.
101.0000000000,5562.8,2505.4,2666.3,25225.
102.0000000000,5562.4,2505.1,2666.2,25225.
103.0000000000,5562.0,2504.8,2666.0,25225.
104.0000000000,5561.6,2504.5,2665.8,25224.
105.0000000000,5561.2,2504.2,2665.6,25224.
106.0000000000,5560.8,2503.9,2665.4,25224.
107.0000000000,5560.3,2503.6,2665.2,25223.
108.0000000000,5559.9,2503.3,2663.4,25223.
109.0000000000,5559.5,2503.0,2663.1,25223.
110.0000000000,5559.1,2502.7,2663.0,25223.
111.0000000000,5558.7,2502.4,2663.0,25222.
112.0000000000,5558.3,2502.2,2663.0,25222.
113.0000000000,5557.9,2501.9,2663.0,25222.
114.0000000000,5557.5,2501.6,2662.9,25222.
115.0000000000,5557.2,2501.4,2662.9,25221.
116.0000000000,5556.8,2501.1,2662.8,25221.
117.0000000000,5556.5,2500.9,2662.6,25221.
118.0000000000,5556.1,2500.7,2657.4,25220.
119.0000000000,5555.8,2500.4,2648.3,25220.
120.0000000000,5555.5,2500.2,2648.2,25220.
121.0000000000,5555.1,2500.0,2649.7,25220.
122.0000000000,5554.8,2499.8,2648.2,25219.
123.0000000000,5554.5,2499.6,2649.7,25219.
124.0000000000,5554.2,2499.4,2651.5,25219.
125.0000000000,5553.9,2499.2,2653.1,25219.
126.0000000000,5553.6,2499.0,2654.5,25218.
127.0000000000,5553.4,2498.8,2655.5,25218.
128.0000000000,5553.1,2498.6,2656.4,25218.
129.0000000000,5552.8,2498.4,2657.1,25218.
130.0000000000,5552.5,2498.2,2655.9,25218.
131.0000000000,5552.3,2498.0,2654.1,25217.
132.0000000000,5552.0,2497.9,2654.4,25217.
133.0000000000,5551.8,2497.7,2655.0,25217.
134.0000000000,5551.5,2497.5,2655.7,25217.
135.0000000000,5551.3,2497.3,2653.5,25216.
136.0000000000,5551.0,2497.2,2653.8,25216.
137.0000000000,5550.8,2497.0,2654.4,25216.
138.0000000000,5550.6,2496.9,2655.0,25216.
139.0000000000,5550.3,2496.7,2655.6,25216.
140.0000000000,5550.1,2496.6,2656.0,25215.
141.0000000000,5549.9,2496.4,2656.3,25215.
142.0000000000,5549.7,2496.3,2656.5,25215.
143.0000000000,5549.4,2496.1,2656.7,25215.
144.0000000000,5549.2,2496.0,2650.7,25215.
145.0000000000,5549.0,2495.9,2649.8,25214.
146.0000000000,5548.8,2495.7,2641.0,25214.
147.0000000000,5548.6,2495.6,2641.3,25214.
148.0000000000,5548.4,2495.5,2643.2,25214.
149.0000000000,5548.2,2495.4,2644.0,25214.
150.0000000000,5548.0,2495.2,2645.8,25213.
151.0000000000,5547.8,2495.1,2647.6,25213.
152.0000000000,5547.7,2495.0,2649.1,25213.
153.0000000000,5547.5,2494.9,2650.4,25213.
154.0000000000,5547.3,2494.7,2651.1,25213.
155.0000000000,5547.1,2494.6,2651.9,25213.
156.0000000000,5547.0,2494.5,2652.5,25212.
157.0000000000,5546.8,2494.4,2653.0,25212.
158.0000000000,5546.6,2494.3,2653.3,25212.
159.0000000000,5546.5,2494.2,2651.4,25212.
160.0000000000,5546.3,2494.0,2651.5,25212.
161.0000000000,5546.2,2493.9,2651.9,25212.
162.0000000000,5546.0,2493.8,2652.3,25212.
163.0000000000,5545.9,2493.7,2652.6,25211.
164.0000000000,5545.7,2493.6,2652.9,25211.
165.0000000000,5545.6,2493.5,2651.8,25211.
166.0000000000,5545.5,2493.4,2639.7,25211.
167.0000000000,5545.3,2493.3,2638.4,25211.
168.0000000000,5545.2,2493.2,2639.9,25211.
169.0000000000,5545.1,2493.1,2641.1,25210.
170.0000000000,5544.9,2493.0,2642.8,25210.
171.0000000000,5544.8,2492.9,2644.7,25210.
172.0000000000,5544.7,2492.8,2646.3,25210.
173.0000000000,5544.6,2492.7,2647.6,25210.
174.0000000000,5544.4,2492.6,2648.7,25210.
175.0000000000,5544.3,2492.5,2649.6,25210.
176.0000000000,5544.2,2492.4,2650.2,25210.
177.0000000000,5544.1,2492.4,2650.8,25209.
178.0000000000,5544.0,2492.3,2651.2,25209.
179.0000000000,5543.9,2492.2,2651.5,25209.
180.0000000000,5543.7,2492.1,2651.7,25209.
181.0000000000,5543.6,2492.0,2648.9,25209.
182.0000000000,5543.5,2491.9,2648.8,25209.
183.0000000000,5543.4,2491.8,2648.5,25209.
184.0000000000,5543.3,2491.7,2649.0,25209.
185.0000000000,5543.2,2491.6,2649.5,25209.
186.0000000000,5543.1,2491.5,2650.0,25209.
187.0000000000,5543.0,2491.5,2650.5,25208.
188.0000000000,5542.9,2491.4,2650.8,25208.
189.0000000000,5542.8,2491.3,2651.1,25208.
190.0000000000,5542.7,2491.2,2651.3,25208.
191.0000000000,5542.6,2491.1,2651.4,25208.
192.0000000000,5542.5,2491.0,2651.5,25208.
193.0000000000,5542.4,2490.9,2651.6,25208.
194.0000000000,5542.3,2490.9,2651.7,25208.
195.0000000000,5542.2,2490.8,2651.7,25208.
196.0000000000,5542.1,2490.7,2651.0,25208.
197.0000000000,5542.0,2490.6,2643.0,25208.
198.0000000000,5541.9,2490.5,2638.4,25207.
199.0000000000,5541.8,2490.4,2638.4,25207.
200.0000000000,5541.7,2490.4,2638.8,25207.
201.0000000000,5541.6,2490.3,2640.6,25207.
202.0000000000,5541.5,2490.2,2642.2,25207.
203.0000000000,5541.4,2490.1,2643.5,25207.
204.0000000000,5541.3,2490.0,2644.9,25207.
205.0000000000,5541.2,2489.9,2646.1,25207.
206.0000000000,5541.2,2489.9,2647.1,25207.
207.0000000000,5541.1,2489.8,2647.9,25207.
208.0000000000,5541.0,2489.7,2648.2,25207.
209.0000000000,5540.9,2489.6,2648.7,25207.
210.0000000000,5540.8,2489.5,2647.9,25206.
211.0000000000,5540.7,2489.5,2648.2,25206.
212.0000000000,5540.6,2489.4,2648.6,25206.
213.0000000000,5540.5,2489.3,2649.0,25206.
214.0000000000,5540.5,2489.2,2649.4,25206.
215.0000000000,5540.4,2489.1,2649.6,25206.
216.0000000000,5540.3,2489.1,2649.9,25206.
217.0000000000,5540.2,2489.0,2650.0,25206.
218.0000000000,5540.1,2488.9,2650.2,25206.
219.0000000000,5540.0,2488.8,2650.3,25206.
220.0000000000,5539.8,2488.7,2650.4,25206.
221.0000000000,5539.6,2488.7,2650.4,25206.
222.0000000000,5539.4,2488.6,2650.5,25206.
223.0000000000,5539.2,2488.5,2650.4,25205.
224.0000000000,5539.1,2488.4,2650.1,25205.
225.0000000000,5539.0,2488.3,2650.1,25205.
226.0000000000,5538.9,2488.3,2650.1,25205.
227.0000000000,5538.7,2488.2,2650.2,25205.
228.0000000000,5538.6,2488.1,2650.2,25205.
229.0000000000,5538.4,2488.0,2650.3,25205.
230.0000000000,5538.3,2488.0,2650.3,25205.
231.0000000000,5538.1,2487.9,2650.4,25205.
232.0000000000,5538.0,2487.8,2650.4,25205.
233.0000000000,5537.9,2487.7,2650.4,25205.
234.0000000000,5537.8,2487.7,2650.1,25205.
235.0000000000,5537.7,2487.6,2650.1,25205.
236.0000000000,5537.6,2487.5,2643.8,25205.
237.0000000000,5537.5,2487.4,2643.3,25204.
238.0000000000,5537.4,2487.3,2643.1,25204.
239.0000000000,5537.3,2487.3,2635.8,25204.
240.0000000000,5537.2,2487.2,2629.7,25204.
241.0000000000,5537.2,2487.1,2631.1,25204.
242.0000000000,5537.1,2487.0,2633.8,25204.
243.0000000000,5537.0,2487.0,2636.6,25204.
244.0000000000,5536.9,2486.9,2639.1,25204.
245.0000000000,5536.8,2486.8,2641.2,25204.
246.0000000000,5536.7,2486.7,2640.0,25204.
247.0000000000,5536.7,2486.7,2641.2,25204.
248.0000000000,5536.6,2486.6,2640.3,25204.
249.0000000000,5536.5,2486.5,2640.1,25204.
250.0000000000,5536.4,2486.4,2641.4,25204.
251.0000000000,5536.3,2486.4,2642.7,25204.
252.0000000000,5536.3,2486.3,2642.1,25203.
253.0000000000,5536.2,2486.2,2642.8,25203.
254.0000000000,5536.1,2486.1,2642.9,25203.
255.0000000000,5536.0,2486.1,2643.8,25203.
256.0000000000,5536.0,2486.0,2644.8,25203.
257.0000000000,5535.9,2485.9,2645.6,25203.
258.0000000000,5535.8,2485.9,2646.3,25203.
259.0000000000,5535.7,2485.8,2646.9,25203.
260.0000000000,5535.7,2485.7,2645.8,25203.
261.0000000000,5535.6,2485.6,2643.0,25203.
262.0000000000,5535.5,2485.6,2642.6,25203.
263.0000000000,5535.5,2485.5,2625.2,25203.
264.0000000000,5535.4,2485.4,2610.4,25203.
265.0000000000,5535.3,2485.4,2612.3,25203.
266.0000000000,5535.2,2485.3,2617.3,25203.
267.0000000000,5535.2,2485.2,2622.6,25203.
268.0000000000,5535.1,2485.1,2627.4,25203.
269.0000000000,5535.0,2485.1,2631.4,25202.
270.0000000000,5535.0,2485.0,2634.7,25202.
271.0000000000,5534.9,2484.9,2637.4,25202.
272.0000000000,5534.8,2484.9,2637.0,25202.
273.0000000000,5534.8,2484.8,2638.6,25202.
274.0000000000,5534.7,2484.7,2640.2,25202.
275.0000000000,5534.6,2484.7,2641.6,25202.
276.0000000000,5534.5,2484.6,2642.8,25202.
277.0000000000,5534.5,2484.5,2643.7,25202.
278.0000000000,5534.4,2484.5,2644.5,25202.
279.0000000000,5534.3,2484.4,2645.1,25202.
280.0000000000,5534.3,2484.3,2645.6,25202.
281.0000000000,5534.2,2484.3,2646.0,25202.
282.0000000000,5534.1,2484.2,2646.3,25202.
283.0000000000,5534.1,2484.2,2646.6,25202.
284.0000000000,5534.0,2484.1,2646.7,25202.
285.0000000000,5534.0,2484.0,2646.9,25202.
286.0000000000,5533.9,2484.0,2647.0,25202.
287.0000000000,5533.8,2483.9,2644.8,25202.
288.0000000000,5533.8,2483.8,2640.8,25202.
289.0000000000,5533.7,2483.8,2628.6,25202.
290.0000000000,5533.6,2483.7,2628.4,25201.
291.0000000000,5533.6,2483.6,2630.7,25201.
292.0000000000,5533.5,2483.6,2633.3,25201.
293.0000000000,5533.5,2483.5,2635.8,25201.
294.0000000000,5533.4,2483.5,2638.0,25201.
295.0000000000,5533.3,2483.4,2639.8,25201.
296.0000000000,5533.3,2483.3,2641.3,25201.
297.0000000000,5533.2,2483.3,2642.4,25201.
298.0000000000,5533.2,2483.2,2643.4,25201.
299.0000000000,5533.1,2483.2,2644.1,25201.
300.0000000000,5533.0,2483.1,2644.7,25201.
301.0000000000,5533.0,2483.0,2645.2,25201.
302.0000000000,5532.9,2483.0,2645.6,25201.
303.0000000000,5532.9,2482.9,2645.9,25201.
304.0000000000,5532.8,2482.9,2646.0,25201.
305.0000000000,5532.8,2482.8,2646.2,25201.
306.0000000000,5532.7,2482.8,2646.4,25201.
307.0000000000,5532.6,2482.7,2646.5,25201.
308.0000000000,5532.6,2482.7,2645.1,25201.
309.0000000000,5532.5,2482.6,2644.6,25201.
310.0000000000,5532.5,2482.6,2643.5,25201.
311.0000000000,5532.4,2482.5,2642.7,25201.
312.0000000000,5532.4,2482.5,2643.1,25201.
313.0000000000,5532.3,2482.5,2642.5,25201.
314.0000000000,5532.3,2482.4,2643.0,25201.
315.0000000000,5532.3,2482.4,2643.7,25201.
316.0000000000,5532.2,2482.3,2644.0,25200.
317.0000000000,5532.2,2482.3,2644.5,25200.
318.0000000000,5532.1,2482.2,2645.0,25200.
319.0000000000,5532.1,2482.2,2645.4,25200.
320.0000000000,5532.0,2482.2,2645.8,25200.
321.0000000000,5532.0,2482.1,2646.1,25200.
322.0000000000,5532.0,2482.1,2646.4,25200.
323.0000000000,5531.9,2482.1,2646.6,25200.
324.0000000000,5531.9,2482.0,2646.7,25200.
325.0000000000,5531.8,2482.0,2646.9,25200.
326.0000000000,5531.8,2482.0,2646.5,25200.
327.0000000000,5531.8,2481.9,2646.1,25200.
328.0000000000,5531.7,2481.9,2642.9,25200.
329.0000000000,5531.7,2481.9,2640.3,25200.
330.0000000000,5531.7,2481.8,2640.6,25200.
331.0000000000,5531.6,2481.8,2641.6,25200.
332.0000000000,5531.6,2481.8,2642.6,25200.
333.0000000000,5531.6,2481.8,2643.5,25200.
334.0000000000,5531.5,2481.7,2644.3,25200.
335.0000000000,5531.5,2481.7,2644.9,25200.
336.0000000000,5531.5,2481.7,2645.5,25200.
337.0000000000,5531.4,2481.7,2645.9,25200.
338.0000000000,5531.4,2481.6,2646.3,25200.
339.0000000000,5531.4,2481.6,2646.6,25200.
340.0000000000,5531.3,2481.6,2646.2,25200.
341.0000000000,5531.3,2481.6,2646.3,25200.
342.0000000000,5531.3,2481.5,2646.6,25200.
343.0000000000,5531.3,2481.5,2646.8,25200.
344.0000000000,5531.2,2481.5,2647.0,25200.
345.0000000000,5531.2,2481.5,2647.2,25200.
346.0000000000,5531.2,2481.4,2647.3,25200.
347.0000000000,5531.2,2481.4,2647.5,25200.
348.0000000000,5531.1,2481.4,2647.6,25200.
349.0000000000,5531.1,2481.4,2647.7,25200.
350.0000000000,5531.1,2481.4,2647.8,25200.
351.0000000000,5531.1,2481.4,2647.9,25200.
352.0000000000,5531.0,2481.3,2647.9,25200.
353.0000000000,5531.0,2481.3,2648.0,25200.
354.0000000000,5531.0,2481.3,2648.1,25200.
355.0000000000,5531.0,2481.3,2645.7,25200.
356.0000000000,5531.0,2481.3,2644.7,25200.
357.0000000000,5530.9,2481.2,2645.0,25200.
358.0000000000,5530.9,2481.2,2645.5,25200.
359.0000000000,5530.9,2481.2,2646.0,25200.
360.0000000000,5530.9,2481.2,2645.6,25200.
361.0000000000,5530.9,2481.2,2644.4,25200.
362.0000000000,5530.8,2481.2,2643.3,25200.
363.0000000000,5530.8,2481.2,2643.8,25200.
364.0000000000,5530.8,2481.1,2644.5,25199.
365.0000000000,5530.8,2481.1,2645.3,25199.
366.0000000000,5530.8,2481.1,2645.9,25199.
367.0000000000,5530.8,2481.1,2646.5,25199.
368.0000000000,5530.8,2481.1,2646.9,25199.
369.0000000000,5530.7,2481.1,2647.3,25199.
370.0000000000,5530.7,2481.1,2647.6,25199.
371.0000000000,5530.7,2481.0,2647.9,25199.
372.0000000000,5530.7,2481.0,2648.1,25199.
373.0000000000,5530.7,2481.0,2648.3,25199.
374.0000000000,5530.7,2481.0,2648.4,25199.
375.0000000000,5530.7,2481.0,2648.6,25199.
376.0000000000,5530.7,2481.0,2648.7,25199.
377.0000000000,5530.6,2481.0,2648.8,25199.
378.0000000000,5530.6,2481.0,2648.9,25199.
379.0000000000,5530.6,2481.0,2649.0,25199.
380.0000000000,5530.6,2481.0,2649.1,25199.
381.0000000000,5530.6,2480.9,2649.1,25199.
382.0000000000,5530.6,2480.9,2649.2,25199.
383.0000000000,5530.6,2480.9,2649.3,25199.
384.0000000000,5530.6,2480.9,2649.3,25199.
385.0000000000,5530.6,2480.9,2649.4,25199.
386.0000000000,5530.6,2480.9,2649.4,25199.
387.0000000000,5530.5,2480.9,2649.5,25199.
388.0000000000,5530.5,2480.9,2649.6,25199.
389.0000000000,5530.5,2480.9,2649.4,25199.
390.0000000000,5530.5,2480.9,2649.4,25199.
391.0000000000,5530.5,2480.9,2649.5,25199.
392.0000000000,5530.5,2480.9,2649.5,25199.
393.0000000000,5530.5,2480.9,2649.6,25199.
394.0000000000,5530.5,2480.9,2649.7,25199.
395.0000000000,5530.5,2480.9,2649.8,25199.
396.0000000000,5530.5,2480.9,2649.8,25199.
397.0000000000,5530.4,2480.8,2649.9,25199.
398.0000000000,5530.4,2480.8,2649.9,25199.
399.0000000000,5530.4,2480.8,2650.0,25199.
400.0000000000,5530.4,2480.8,2650.1,25199.
401.0000000000,5530.4,2480.8,2650.1,25199.
402.0000000000,5530.4,2480.8,2650.2,25199.
403.0000000000,5530.4,2480.8,2650.2,25199.
404.0000000000,5530.4,2480.8,2650.3,25199.
405.0000000000,5530.4,2480.8,2650.4,25199.
406.0000000000,5530.4,2480.8,2650.4,25199.
407.0000000000,5530.4,2480.8,2650.5,25199.
408.0000000000,5530.4,2480.8,2650.5,25200.
409.0000000000,5530.4,2480.8,2650.6,25200.
410.0000000000,5530.3,2480.8,2650.7,25200.
411.0000000000,5530.3,2480.8,2650.7,25200.
412.0000000000,5530.3,2480.8,2650.8,25200.
413.0000000000,5530.3,2480.8,2650.9,25200.
414.0000000000,5530.3,2480.8,2650.9,25200.
415.0000000000,5530.3,2480.8,2651.0,25200.
416.0000000000,5530.3,2480.8,2651.0,25200.
417.0000000000,5530.3,2480.8,2651.1,25200.
418.0000000000,5530.3,2480.8,2651.2,25200.
419.0000000000,5530.3,2480.8,2651.2,25200.
420.0000000000,5530.3,2480.8,2651.3,25200.
421.0000000000,5530.3,2480.8,2651.2,25200.
422.0000000000,5530.3,2480.8,2649.2,25200.
423.0000000000,5530.3,2480.8,2648.5,25200.
424.0000000000,5530.3,2480.8,2648.7,25200.
425.0000000000,5530.3,2480.8,2649.2,25200.
426.0000000000,5530.3,2480.8,2649.6,25200.
427.0000000000,5530.3,2480.8,2650.0,25200.
428.0000000000,5530.3,2480.8,2650.4,25200.
429.0000000000,5530.4,2480.8,2650.7,25200.
430.0000000000,5530.4,2480.8,2651.0,25200.
431.0000000000,5530.4,2480.8,2651.2,25200.
432.0000000000,5530.4,2480.8,2651.4,25200.
433.0000000000,5530.4,2480.8,2651.6,25200.
434.0000000000,5530.4,2480.8,2651.7,25200.
435.0000000000,5530.4,2480.8,2651.8,25200.
436.0000000000,5530.4,2480.8,2651.9,25200.
437.0000000000,5530.4,2480.8,2652.0,25200.
438.0000000000,5530.4,2480.8,2652.1,25200.
439.0000000000,5530.4,2480.8,2652.2,25200.
440.0000000000,5530.4,2480.8,2652.3,25200.
441.0000000000,5530.5,2480.8,2652.4,25200.
442.0000000000,5530.5,2480.8,2652.5,25200.
443.0000000000,5530.5,2480.8,2652.6,25200.
444.0000000000,5530.5,2480.8,2652.7,25200.
445.0000000000,5530.5,2480.8,2652.8,25200.
446.0000000000,5530.5,2480.8,2652.8,25200.
447.0000000000,5530.5,2480.8,2652.9,25200.
448.0000000000,5530.6,2480.8,2652.5,25200.
449.0000000000,5530.6,2480.8,2652.5,25200.
450.0000000000,5530.6,2480.8,2652.7,25200.
451.0000000000,5530.6,2480.8,2652.7,25200.
452.0000000000,5530.6,2480.8,2652.9,25200.
453.0000000000,5530.6,2480.8,2653.0,25200.
454.0000000000,5530.7,2480.8,2653.1,25200.
455.0000000000,5530.7,2480.8,2653.3,25200.
456.0000000000,5530.7,2480.8,2653.4,25200.
457.0000000000,5530.7,2480.8,2653.5,25200.
458.0000000000,5530.7,2480.8,2653.6,25200.
459.0000000000,5530.8,2480.8,2651.9,25200.
460.0000000000,5530.8,2480.8,2651.9,25201.
461.0000000000,5530.8,2480.8,2652.1,25201.
462.0000000000,5530.8,2480.8,2652.4,25201.
463.0000000000,5530.8,2480.8,2652.5,25201.
464.0000000000,5530.9,2480.8,2652.8,25201.
465.0000000000,5530.9,2480.8,2653.1,25201.
466.0000000000,5530.9,2480.8,2653.4,25201.
467.0000000000,5530.9,2480.8,2653.6,25201.
468.0000000000,5530.9,2480.8,2653.8,25201.
469.0000000000,5531.0,2480.8,2654.0,25201.
470.0000000000,5531.0,2480.8,2654.2,25201.
471.0000000000,5531.0,2480.8,2654.3,25201.
472.0000000000,5531.0,2480.8,2654.5,25201.
473.0000000000,5531.1,2480.8,2654.6,25201.
474.0000000000,5531.1,2480.8,2654.7,25201.
475.0000000000,5531.1,2480.8,2654.6,25201.
476.0000000000,5531.1,2480.8,2654.7,25201.
477.0000000000,5531.1,2480.8,2654.8,25201.
478.0000000000,5531.2,2480.8,2654.9,25201.
479.0000000000,5531.2,2480.8,2655.0,25201.
480.0000000000,5531.2,2480.8,2655.1,25201.
481.0000000000,5531.2,2480.9,2655.3,25201.
482.0000000000,5531.3,2480.9,2655.4,25201.
483.0000000000,5531.3,2480.9,2655.5,25201.
484.0000000000,5531.3,2480.9,2655.6,25201.
485.0000000000,5531.3,2480.9,2655.7,25201.
486.0000000000,5531.4,2480.9,2655.7,25201.
487.0000000000,5531.4,2480.9,2655.8,25202.
488.0000000000,5531.4,2480.9,2655.9,25202.
489.0000000000,5531.4,2480.9,2656.0,25202.
490.0000000000,5531.5,2480.9,2656.1,25202.
491.0000000000,5531.5,2480.9,2656.2,25202.
492.0000000000,5531.5,2480.9,2654.9,25202.
493.0000000000,5531.6,2480.9,2654.9,25202.
494.0000000000,5531.6,2480.9,2654.5,25202.
495.0000000000,5531.6,2480.9,2653.6,25202.
496.0000000000,5531.6,2480.9,2653.8,25202.
497.0000000000,5531.7,2480.9,2654.3,25202.
498.0000000000,5531.7,2480.9,2653.4,25202.
499.0000000000,5531.7,2480.9,2653.5,25202.
500.0000000000,5531.8,2480.9,2654.0,25202.
501.0000000000,5531.8,2480.9,2654.6,25202.
502.0000000000,5531.8,2480.9,2655.1,25202.
503.0000000000,5531.8,2480.9,2655.5,25202.
504.0000000000,5531.9,2480.9,2655.9,25202.
505.0000000000,5531.9,2481.0,2656.3,25202.
506.0000000000,5531.9,2481.0,2656.5,25202.
507.0000000000,5532.0,2481.0,2656.8,25203.
508.0000000000,5532.0,2481.0,2656.5,25203.
509.0000000000,5532.0,2481.0,2656.6,25203.
510.0000000000,5532.0,2481.0,2655.5,25203.
511.0000000000,5532.1,2481.0,2647.2,25203.
512.0000000000,5532.1,2481.0,2646.5,25203.
513.0000000000,5532.1,2481.0,2647.7,25203.
514.0000000000,5532.2,2481.0,2649.4,25203.
515.0000000000,5532.2,2481.0,2651.0,25203.
516.0000000000,5532.2,2481.0,2652.4,25203.
517.0000000000,5532.3,2481.0,2653.5,25203.
518.0000000000,5532.3,2481.0,2654.5,25203.
519.0000000000,5532.3,2481.0,2655.3,25203.
520.0000000000,5532.3,2481.0,2656.0,25203.
521.0000000000,5532.4,2481.0,2656.5,25203.
522.0000000000,5532.4,2481.0,2657.0,25203.
523.0000000000,5532.4,2481.0,2657.3,25203.
524.0000000000,5532.5,2481.0,2657.6,25204.
525.0000000000,5532.5,2481.0,2657.8,25204.
526.0000000000,5532.5,2481.0,2657.9,25204.
527.0000000000,5532.6,2481.0,2658.1,25204.
528.0000000000,5532.6,2481.1,2658.0,25204.
529.0000000000,5532.6,2481.1,2656.5,25204.
530.0000000000,5532.7,2481.1,2653.3,25204.
531.0000000000,5532.7,2481.1,2653.5,25204.
532.0000000000,5532.7,2481.1,2654.3,25204.
533.0000000000,5532.8,2481.1,2655.2,25204.
534.0000000000,5532.8,2481.1,2656.0,25204.
535.0000000000,5532.8,2481.1,2656.7,25204.
536.0000000000,5532.9,2481.1,2638.6,25204.
537.0000000000,5532.9,2481.1,2630.2,25204.
538.0000000000,5532.9,2481.1,2629.6,25204.
539.0000000000,5532.9,2481.1,2633.4,25204.
540.0000000000,5533.0,2481.1,2637.6,25205.
541.0000000000,5533.0,2481.1,2634.8,25205.
542.0000000000,5533.0,2481.1,2637.8,25205.
543.0000000000,5533.1,2481.1,2641.5,25205.
544.0000000000,5533.1,2481.1,2644.7,25205.
545.0000000000,5533.1,2481.1,2647.6,25205.
546.0000000000,5533.2,2481.1,2650.0,25205.
547.0000000000,5533.2,2481.1,2651.9,25205.
548.0000000000,5533.2,2481.1,2653.5,25205.
549.0000000000,5533.3,2481.1,2654.7,25205.
550.0000000000,5533.3,2481.1,2655.8,25205.
551.0000000000,5533.3,2481.1,2656.6,25205.
552.0000000000,5533.4,2481.2,2657.3,25205.
553.0000000000,5533.4,2481.2,2657.9,25205.
554.0000000000,5533.4,2481.2,2658.3,25205.
555.0000000000,5533.5,2481.2,2658.7,25206.
556.0000000000,5533.5,2481.2,2658.9,25206.
557.0000000000,5533.5,2481.2,2659.1,25206.
558.0000000000,5533.6,2481.2,2657.9,25206.
559.0000000000,5533.6,2481.2,2658.0,25206.
560.0000000000,5533.6,2481.2,2658.4,25206.
561.0000000000,5533.7,2481.2,2658.8,25206.
562.0000000000,5533.7,2481.2,2657.3,25206.
563.0000000000,5533.7,2481.2,2655.3,25206.
564.0000000000,5533.8,2481.2,2654.0,25206.
565.0000000000,5533.8,2481.2,2654.6,25206.
566.0000000000,5533.8,2481.2,2655.6,25206.
567.0000000000,5533.9,2481.2,2656.6,25206.
568.0000000000,5533.9,2481.2,2657.5,25206.
569.0000000000,5533.9,2481.2,2658.2,25206.
570.0000000000,5534.0,2481.2,2658.8,25207.
571.0000000000,5534.0,2481.2,2658.6,25207.
572.0000000000,5534.0,2481.2,2658.9,25207.
573.0000000000,5534.1,2481.2,2659.4,25207.
574.0000000000,5534.1,2481.2,2659.8,25207.
575.0000000000,5534.2,2481.2,2660.2,25207.
576.0000000000,5534.2,2481.3,2660.5,25207.
577.0000000000,5534.2,2481.3,2660.8,25207.
578.0000000000,5534.3,2481.3,2661.0,25207.
579.0000000000,5534.3,2481.3,2657.9,25207.
580.0000000000,5534.3,2481.3,2649.3,25207.
581.0000000000,5534.4,2481.3,2649.3,25207.
582.0000000000,5534.4,2481.3,2650.8,25207.
583.0000000000,5534.4,2481.3,2652.7,25208.
584.0000000000,5534.5,2481.3,2654.5,25208.
585.0000000000,5534.5,2481.3,2656.0,25208.
586.0000000000,5534.6,2481.3,2657.2,25208.
587.0000000000,5534.6,2481.3,2658.3,25208.
588.0000000000,5534.6,2481.3,2659.2,25208.
589.0000000000,5534.7,2481.3,2659.0,25208.
590.0000000000,5534.7,2481.3,2657.4,25208.
591.0000000000,5534.7,2481.3,2657.8,25208.
592.0000000000,5534.8,2481.3,2658.6,25208.
593.0000000000,5534.8,2481.3,2659.4,25208.
594.0000000000,5534.8,2481.3,2659.5,25208.
595.0000000000,5534.9,2481.3,2657.4,25208.
596.0000000000,5534.9,2481.3,2654.5,25208.
597.0000000000,5535.0,2481.3,2655.1,25209.
598.0000000000,5535.0,2481.3,2656.3,25209.
599.0000000000,5535.0,2481.3,2657.5,25209.
600.0000000000,5535.1,2481.3,2658.6,25209.
601.0000000000,5535.1,2481.4,2659.5,25209.
602.0000000000,5535.1,2481.4,2660.3,25209.
603.0000000000,5535.2,2481.4,2661.0,25209.
604.0000000000,5535.2,2481.4,2661.5,25209.
605.0000000000,5535.2,2481.4,2661.9,25209.
606.0000000000,5535.3,2481.4,2662.3,25209.
607.0000000000,5535.3,2481.4,2662.2,25209.
608.0000000000,5535.4,2481.4,2662.4,25209.
609.0000000000,5535.4,2481.4,2662.6,25209.
610.0000000000,5535.4,2481.4,2662.9,25210.
611.0000000000,5535.5,2481.4,2663.2,25210.
612.0000000000,5535.5,2481.4,2663.4,25210.
613.0000000000,5535.5,2481.4,2660.9,25210.
614.0000000000,5535.6,2481.4,2660.2,25210.
615.0000000000,5535.6,2481.4,2660.6,25210.
616.0000000000,5535.6,2481.4,2659.2,25210.
617.0000000000,5535.7,2481.4,2659.7,25210.
618.0000000000,5535.7,2481.4,2660.5,25210.
619.0000000000,5535.8,2481.4,2661.3,25210.
620.0000000000,5535.8,2481.4,2661.9,25210.
621.0000000000,5535.8,2481.4,2661.7,25210.
622.0000000000,5535.9,2481.4,2661.6,25210.
623.0000000000,5535.9,2481.4,2662.0,25211.
624.0000000000,5535.9,2481.4,2662.6,25211.
625.0000000000,5536.0,2481.4,2662.6,25211.
626.0000000000,5536.0,2481.4,2663.0,25211.
627.0000000000,5536.0,2481.4,2658.9,25211.
628.0000000000,5536.1,2481.5,2658.6,25211.
629.0000000000,5536.1,2481.5,2657.1,25211.
630.0000000000,5536.2,2481.5,2656.7,25211.
631.0000000000,5536.2,2481.5,2657.8,25211.
632.0000000000,5536.2,2481.5,2659.1,25211.
633.0000000000,5536.3,2481.5,2660.3,25211.
634.0000000000,5536.3,2481.5,2661.3,25211.
635.0000000000,5536.3,2481.5,2652.1,25211.
636.0000000000,5536.4,2481.5,2650.5,25212.
637.0000000000,5536.4,2481.5,2652.1,25212.
638.0000000000,5536.4,2481.5,2654.3,25212.
639.0000000000,5536.5,2481.5,2656.4,25212.
640.0000000000,5536.5,2481.5,2658.3,25212.
641.0000000000,5536.6,2481.5,2659.8,25212.
642.0000000000,5536.6,2481.5,2661.1,25212.
643.0000000000,5536.6,2481.5,2662.2,25212.
644.0000000000,5536.7,2481.5,2663.0,25212.
645.0000000000,5536.7,2481.5,2663.7,25212.
646.0000000000,5536.7,2481.5,2664.3,25212.
647.0000000000,5536.8,2481.5,2664.8,25212.
648.0000000000,5536.8,2481.5,2665.2,25212.
649.0000000000,5536.8,2481.5,2661.3,25213.
650.0000000000,5536.9,2481.5,2661.4,25213.
651.0000000000,5536.9,2481.5,2662.0,25213.
652.0000000000,5537.0,2481.5,2662.9,25213.
653.0000000000,5537.0,2481.5,2663.6,25213.
654.0000000000,5537.0,2481.5,2664.3,25213.
655.0000000000,5537.1,2481.5,2664.9,25213.
656.0000000000,5537.1,2481.5,2665.4,25213.
657.0000000000,5537.1,2481.5,2665.8,25213.
658.0000000000,5537.2,2481.5,2666.1,25213.
659.0000000000,5537.2,2481.5,2666.2,25213.
660.0000000000,5537.2,2481.5,2665.7,25213.
661.0000000000,5537.3,2481.5,2663.5,25214.
662.0000000000,5537.3,2481.5,2663.6,25214.
663.0000000000,5537.3,2481.5,2664.2,25214.
664.0000000000,5537.4,2481.6,2664.8,25214.
665.0000000000,5537.4,2481.6,2665.4,25214.
666.0000000000,5537.4,2481.6,2665.9,25214.
667.0000000000,5537.5,2481.6,2666.4,25214.
668.0000000000,5537.5,2481.6,2666.8,25214.
669.0000000000,5537.6,2481.6,2667.1,25214.
670.0000000000,5537.6,2481.6,2667.4,25214.
671.0000000000,5537.6,2481.6,2667.6,25214.
672.0000000000,5537.7,2481.6,2667.8,25214.
673.0000000000,5537.7,2481.6,2668.0,25215.
674.0000000000,5537.7,2481.6,2654.1,25215.
675.0000000000,5537.8,2481.6,2645.7,25215.
676.0000000000,5537.8,2481.6,2646.7,25215.
677.0000000000,5537.8,2481.6,2649.5,25215.
678.0000000000,5537.9,2481.6,2652.7,25215.
679.0000000000,5537.9,2481.6,2655.7,25215.
680.0000000000,5537.9,2481.6,2658.2,25215.
681.0000000000,5538.0,2481.6,2660.3,25215.
682.0000000000,5538.0,2481.6,2662.1,25215.
683.0000000000,5538.0,2481.6,2663.5,25215.
684.0000000000,5538.1,2481.6,2664.6,25215.
685.0000000000,5538.1,2481.6,2665.5,25216.
686.0000000000,5538.2,2481.6,2666.3,25216.
687.0000000000,5538.2,2481.6,2666.9,25216.
688.0000000000,5538.2,2481.6,2667.4,25216.
689.0000000000,5538.3,2481.6,2667.8,25216.
690.0000000000,5538.3,2481.6,2668.2,25216.
691.0000000000,5538.3,2481.6,2668.4,25216.
692.0000000000,5538.4,2481.6,2667.4,25216.
693.0000000000,5538.4,2481.6,2667.6,25216.
694.0000000000,5538.4,2481.6,2667.9,25216.
695.0000000000,5538.5,2481.6,2668.2,25216.
696.0000000000,5538.5,2481.6,2668.6,25216.
697.0000000000,5538.5,2481.6,2668.9,25217.
698.0000000000,5538.6,2481.6,2669.1,25217.
699.0000000000,5538.6,2481.6,2669.4,25217.
700.0000000000,5538.6,2481.6,2669.6,25217.
701.0000000000,5538.7,2481.6,2669.7,25217.
702.0000000000,5538.7,2481.6,2669.9,25217.
703.0000000000,5538.7,2481.6,2670.0,25217.
704.0000000000,5538.8,2481.6,2670.2,25217.
705.0000000000,5538.8,2481.6,2670.3,25217.
706.0000000000,5538.8,2481.6,2670.4,25217.
707.0000000000,5538.9,2481.6,2670.5,25217.
708.0000000000,5538.9,2481.6,2670.6,25217.
709.0000000000,5538.9,2481.6,2670.7,25218.
710.0000000000,5539.0,2481.6,2670.8,25218.
711.0000000000,5539.0,2481.6,2670.9,25218.
712.0000000000,5539.0,2481.6,2671.0,25218.
713.0000000000,5539.1,2481.6,2671.1,25218.
714.0000000000,5539.1,2481.6,2671.2,25218.
715.0000000000,5539.1,2481.6,2671.3,25218.
716.0000000000,5539.2,2481.6,2671.4,25218.
717.0000000000,5539.2,2481.6,2671.5,25218.
718.0000000000,5539.2,2481.6,2671.4,25218.
719.0000000000,5539.3,2481.6,2671.5,25218.
720.0000000000,5539.3,2481.6,2671.6,25218.
721.0000000000,5539.3,2481.6,2671.7,25219.
722.0000000000,5539.4,2481.6,2671.7,25219.
723.0000000000,5539.4,2481.6,2671.6,25219.
724.0000000000,5539.4,2481.6,2671.8,25219.
725.0000000000,5539.5,2481.6,2671.9,25219.
726.0000000000,5539.5,2481.6,2672.0,25219.
727.0000000000,5539.5,2481.6,2666.8,25219.
728.0000000000,5539.6,2481.6,2666.3,25219.
729.0000000000,5539.6,2481.6,2667.0,25219.
730.0000000000,5539.6,2481.6,2667.6,25219.
731.0000000000,5539.7,2481.6,2667.5,25219.
732.0000000000,5539.7,2481.6,2666.6,25220.
733.0000000000,5539.7,2481.6,2665.5,25220.
734.0000000000,5539.8,2481.6,2666.3,25220.
735.0000000000,5539.8,2481.6,2667.5,25220.
736.0000000000,5539.8,2481.6,2668.5,25220.
737.0000000000,5539.9,2481.6,2669.5,25220.
738.0000000000,5539.9,2481.6,2670.2,25220.
739.0000000000,5539.9,2481.6,2670.8,25220.
740.0000000000,5540.0,2481.6,2668.7,25220.
741.0000000000,5540.0,2481.6,2668.7,25220.
742.0000000000,5540.0,2481.6,2669.4,25220.
743.0000000000,5540.1,2481.6,2670.1,25220.
744.0000000000,5540.1,2481.6,2670.8,25221.
745.0000000000,5540.1,2481.6,2671.5,25221.
746.0000000000,5540.1,2481.6,2672.0,25221.
747.0000000000,5540.2,2481.6,2672.4,25221.
748.0000000000,5540.2,2481.6,2672.8,25221.
749.0000000000,5540.2,2481.6,2673.1,25221.
750.0000000000,5540.3,2481.6,2673.4,25221.
751.0000000000,5540.3,2481.6,2673.6,25221.
752.0000000000,5540.3,2481.6,2672.0,25221.
753.0000000000,5540.4,2481.6,2670.1,25221.
754.0000000000,5540.4,2481.6,2670.2,25221.
755.0000000000,5540.4,2481.6,2670.8,25222.
756.0000000000,5540.5,2481.6,2671.5,25222.
757.0000000000,5540.5,2481.6,2672.1,25222.
758.0000000000,5540.5,2481.6,2672.7,25222.
759.0000000000,5540.6,2481.6,2673.2,25222.
760.0000000000,5540.6,2481.6,2673.6,25222.
761.0000000000,5540.6,2481.6,2672.3,25222.
762.0000000000,5540.6,2481.6,2670.3,25222.
763.0000000000,5540.7,2481.6,2670.6,25222.
764.0000000000,5540.7,2481.5,2671.3,25222.
765.0000000000,5540.7,2481.5,2671.9,25222.
766.0000000000,5540.8,2481.5,2672.6,25222.
767.0000000000,5540.8,2481.5,2673.2,25223.
768.0000000000,5540.8,2481.5,2673.7,25223.
769.0000000000,5540.9,2481.5,2674.1,25223.
770.0000000000,5540.9,2481.5,2674.5,25223.
771.0000000000,5540.9,2481.5,2674.8,25223.
772.0000000000,5541.0,2481.5,2675.1,25223.
773.0000000000,5541.0,2481.5,2675.3,25223.
774.0000000000,5541.0,2481.5,2675.5,25223.
775.0000000000,5541.0,2481.5,2675.7,25223.
776.0000000000,5541.1,2481.5,2675.9,25223.
777.0000000000,5541.1,2481.5,2676.0,25223.
778.0000000000,5541.1,2481.5,2675.9,25224.
779.0000000000,5541.2,2481.5,2676.0,25224.
780.0000000000,5541.2,2481.5,2676.2,25224.
781.0000000000,5541.2,2481.5,2676.3,25224.
782.0000000000,5541.3,2481.5,2676.5,25224.
783.0000000000,5541.3,2481.5,2676.6,25224.
784.0000000000,5541.3,2481.5,2676.7,25224.
785.0000000000,5541.3,2481.5,2676.8,25224.
786.0000000000,5541.4,2481.5,2676.9,25224.
787.0000000000,5541.4,2481.5,2677.0,25224.
788.0000000000,5541.4,2481.5,2677.1,25224.
789.0000000000,5541.5,2481.4,2676.6,25224.
790.0000000000,5541.5,2481.4,2676.5,25225.
791.0000000000,5541.5,2481.4,2676.5,25225.
792.0000000000,5541.5,2481.4,2676.7,25225.
793.0000000000,5541.6,2481.4,2677.0,25225.
794.0000000000,5541.6,2481.4,2674.8,25225.
795.0000000000,5541.6,2481.4,2674.8,25225.
796.0000000000,5541.7,2481.4,2675.2,25225.
797.0000000000,5541.7,2481.4,2675.0,25225.
798.0000000000,5541.7,2481.4,2675.2,25225.
799.0000000000,5541.8,2481.4,2675.4,25225.
800.0000000000,5541.8,2481.4,2675.9,25225.
801.0000000000,5541.8,2481.4,2676.4,25226.
802.0000000000,5541.8,2481.4,2676.8,25226.
803.0000000000,5541.9,2481.4,2677.2,25226.
804.0000000000,5541.9,2481.4,2677.5,25226.
805.0000000000,5541.9,2481.4,2677.8,25226.
806.0000000000,5542.0,2481.4,2678.1,25226.
807.0000000000,5542.0,2481.4,2677.8,25226.
808.0000000000,5542.0,2481.4,2677.9,25226.
809.0000000000,5542.0,2481.4,2675.4,25226.
810.0000000000,5542.1,2481.4,2665.7,25226.
811.0000000000,5542.1,2481.3,2660.1,25226.
812.0000000000,5542.1,2481.3,2661.4,25227.
813.0000000000,5542.2,2481.3,2664.0,25227.
814.0000000000,5542.2,2481.3,2666.7,25227.
815.0000000000,5542.2,2481.3,2668.7,25227.
816.0000000000,5542.3,2481.3,2670.7,25227.
817.0000000000,5542.3,2481.3,2672.5,25227.
818.0000000000,5542.3,2481.3,2673.9,25227.
819.0000000000,5542.3,2481.3,2675.1,25227.
820.0000000000,5542.4,2481.3,2676.0,25227.
821.0000000000,5542.4,2481.3,2676.8,25227.
822.0000000000,5542.4,2481.3,2677.4,25227.
823.0000000000,5542.5,2481.3,2677.9,25227.
824.0000000000,5542.5,2481.3,2678.4,25228.
825.0000000000,5542.5,2481.3,2678.7,25228.
826.0000000000,5542.5,2481.3,2678.5,25228.
827.0000000000,5542.6,2481.3,2678.8,25228.
828.0000000000,5542.6,2481.3,2678.9,25228.
829.0000000000,5542.6,2481.3,2678.0,25228.
830.0000000000,5542.7,2481.3,2678.2,25228.
831.0000000000,5542.7,2481.3,2678.6,25228.
832.0000000000,5542.7,2481.2,2678.1,25228.
833.0000000000,5542.7,2481.2,2674.2,25228.
834.0000000000,5542.8,2481.2,2674.3,25228.
835.0000000000,5542.8,2481.2,2675.1,25229.
836.0000000000,5542.8,2481.2,2673.9,25229.
837.0000000000,5542.9,2481.2,2674.1,25229.
838.0000000000,5542.9,2481.2,2671.8,25229.
839.0000000000,5542.9,2481.2,2672.6,25229.
840.0000000000,5542.9,2481.2,2673.9,25229.
841.0000000000,5543.0,2481.2,2675.2,25229.
842.0000000000,5543.0,2481.2,2676.3,25229.
843.0000000000,5543.0,2481.2,2677.3,25229.
844.0000000000,5543.1,2481.2,2675.7,25229.
845.0000000000,5543.1,2481.2,2676.2,25229.
846.0000000000,5543.1,2481.2,2677.1,25230.
847.0000000000,5543.1,2481.2,2673.8,25230.
848.0000000000,5543.2,2481.2,2674.3,25230.
849.0000000000,5543.2,2481.2,2675.4,25230.
850.0000000000,5543.2,2481.2,2676.5,25230.
851.0000000000,5543.3,2481.2,2677.5,25230.
852.0000000000,5543.3,2481.2,2678.4,25230.
853.0000000000,5543.3,2481.2,2679.1,25230.
854.0000000000,5543.4,2481.2,2679.7,25230.
855.0000000000,5543.4,2481.1,2680.2,25230.
856.0000000000,5543.4,2481.1,2680.6,25230.
857.0000000000,5543.4,2481.1,2680.8,25231.
858.0000000000,5543.5,2481.1,2681.1,25231.
859.0000000000,5543.5,2481.1,2681.4,25231.
860.0000000000,5543.5,2481.1,2681.6,25231.
861.0000000000,5543.6,2481.1,2669.2,25231.
862.0000000000,5543.6,2481.1,2659.4,25231.
863.0000000000,5543.6,2481.1,2653.6,25231.
864.0000000000,5543.6,2481.1,2653.6,25231.
865.0000000000,5543.7,2481.1,2656.0,25231.
866.0000000000,5543.7,2481.1,2654.9,25231.
867.0000000000,5543.7,2481.1,2649.3,25231.
868.0000000000,5543.8,2481.1,2652.9,25231.
869.0000000000,5543.8,2481.1,2657.5,25232.
870.0000000000,5543.8,2481.1,2662.0,25232.
871.0000000000,5543.8,2481.1,2661.8,25232.
872.0000000000,5543.9,2481.1,2663.9,25232.
873.0000000000,5543.9,2481.1,2666.8,25232.
874.0000000000,5543.9,2481.1,2667.1,25232.
875.0000000000,5544.0,2481.1,2669.2,25232.
876.0000000000,5544.0,2481.1,2670.5,25232.
877.0000000000,5544.0,2481.1,2672.5,25232.
878.0000000000,5544.1,2481.0,2674.3,25232.
879.0000000000,5544.1,2481.0,2665.3,25232.
880.0000000000,5544.1,2481.0,2665.8,25233.
881.0000000000,5544.1,2481.0,2659.8,25233.
882.0000000000,5544.2,2481.0,2661.8,25233.
883.0000000000,5544.2,2481.0,2664.9,25233.
884.0000000000,5544.2,2481.0,2668.0,25233.
885.0000000000,5544.3,2481.0,2670.7,25233.
886.0000000000,5544.3,2481.0,2673.0,25233.
887.0000000000,5544.3,2481.0,2674.9,25233.
888.0000000000,5544.3,2481.0,2676.4,25233.
889.0000000000,5544.4,2481.0,2677.7,25233.
890.0000000000,5544.4,2481.0,2678.7,25233.
891.0000000000,5544.4,2481.0,2679.5,25233.
892.0000000000,5544.5,2481.0,2680.2,25234.
893.0000000000,5544.5,2481.0,2680.7,25234.
894.0000000000,5544.5,2481.0,2680.3,25234.
895.0000000000,5544.5,2481.0,2673.6,25234.
896.0000000000,5544.6,2481.0,2672.9,25234.
897.0000000000,5544.6,2481.0,2670.6,25234.
898.0000000000,5544.6,2481.0,2670.5,25234.
899.0000000000,5544.7,2481.0,2672.0,25234.
900.0000000000,5544.7,2481.0,2673.7,25234.
901.0000000000,5544.7,2481.0,2672.2,25234.
902.0000000000,5544.7,2481.0,2673.2,25234.
903.0000000000,5544.8,2480.9,2674.7,25235.
904.0000000000,5544.8,2480.9,2675.5,25235.
905.0000000000,5544.8,2480.9,2676.7,25235.
906.0000000000,5544.8,2480.9,2677.9,25235.
907.0000000000,5544.9,2480.9,2679.0,25235.
908.0000000000,5544.9,2480.9,2675.7,25235.
909.0000000000,5544.9,2480.9,2672.5,25235.
910.0000000000,5545.0,2480.9,2673.1,25235.
911.0000000000,5545.0,2480.9,2674.6,25235.
912.0000000000,5545.0,2480.9,2675.2,25235.
913.0000000000,5545.0,2480.9,2676.5,25235.
914.0000000000,5545.1,2480.9,2677.8,25236.
915.0000000000,5545.1,2480.9,2679.0,25236.
916.0000000000,5545.1,2480.9,2680.0,25236.
917.0000000000,5545.2,2480.9,2680.8,25236.
918.0000000000,5545.2,2480.9,2681.4,25236.
919.0000000000,5545.2,2480.9,2677.7,25236.
920.0000000000,5545.2,2480.9,2677.9,25236.
921.0000000000,5545.3,2480.9,2678.7,25236.
922.0000000000,5545.3,2480.9,2679.7,25236.
923.0000000000,5545.3,2480.9,2680.5,25236.
924.0000000000,5545.4,2480.9,2681.3,25236.
925.0000000000,5545.4,2480.9,2681.9,25236.
926.0000000000,5545.4,2480.9,2682.5,25237.
927.0000000000,5545.4,2480.9,2682.9,25237.
928.0000000000,5545.5,2480.9,2683.3,25237.
929.0000000000,5545.5,2480.9,2683.6,25237.
930.0000000000,5545.5,2480.9,2683.9,25237.
931.0000000000,5545.5,2480.9,2684.1,25237.
932.0000000000,5545.6,2480.9,2684.3,25237.
933.0000000000,5545.6,2480.9,2684.5,25237.
934.0000000000,5545.6,2480.8,2684.6,25237.
935.0000000000,5545.7,2480.8,2684.8,25237.
936.0000000000,5545.7,2480.8,2684.9,25237.
937.0000000000,5545.7,2480.8,2685.0,25238.
938.0000000000,5545.7,2480.8,2685.1,25238.
939.0000000000,5545.8,2480.8,2685.2,25238.
940.0000000000,5545.8,2480.8,2685.3,25238.
941.0000000000,5545.8,2480.8,2685.4,25238.
942.0000000000,5545.9,2480.8,2685.5,25238.
943.0000000000,5545.9,2480.8,2684.5,25238.
944.0000000000,5545.9,2480.8,2683.3,25238.
945.0000000000,5546.0,2480.8,2683.4,25238.
946.0000000000,5546.0,2480.8,2683.8,25238.
947.0000000000,5546.0,2480.8,2684.2,25238.
948.0000000000,5546.0,2480.8,2684.6,25239.
949.0000000000,5546.1,2480.8,2685.0,25239.
950.0000000000,5546.1,2480.8,2685.3,25239.
951.0000000000,5546.1,2480.8,2685.6,25239.
952.0000000000,5546.1,2480.8,2685.8,25239.
953.0000000000,5546.2,2480.8,2686.0,25239.
954.0000000000,5546.2,2480.8,2686.2,25239.
955.0000000000,5546.2,2480.8,2685.2,25239.
956.0000000000,5546.3,2480.8,2684.3,25239.
957.0000000000,5546.3,2480.8,2682.7,25239.
958.0000000000,5546.3,2480.8,2680.4,25239.
959.0000000000,5546.3,2480.8,2680.9,25240.
960.0000000000,5546.4,2480.8,2681.8,25240.
961.0000000000,5546.4,2480.8,2682.8,25240.
962.0000000000,5546.4,2480.8,2680.1,25240.
963.0000000000,5546.5,2480.8,2679.0,25240.
964.0000000000,5546.5,2480.8,2680.0,25240.
965.0000000000,5546.5,2480.8,2681.2,25240.
966.0000000000,5546.5,2480.8,2682.4,25240.
967.0000000000,5546.6,2480.8,2683.4,25240.
968.0000000000,5546.6,2480.8,2683.6,25240.
969.0000000000,5546.6,2480.8,2683.4,25240.
970.0000000000,5546.7,2480.8,2684.0,25240.
971.0000000000,5546.7,2480.8,2684.7,25241.
972.0000000000,5546.7,2480.8,2685.3,25241.
973.0000000000,5546.8,2480.8,2685.4,25241.
974.0000000000,5546.8,2480.8,2685.9,25241.
975.0000000000,5546.8,2480.8,2686.3,25241.
976.0000000000,5546.9,2480.8,2686.7,25241.
977.0000000000,5546.9,2480.8,2687.1,25241.
978.0000000000,5546.9,2480.8,2687.4,25241.
979.0000000000,5546.9,2480.8,2687.6,25241.
980.0000000000,5547.0,2480.8,2687.9,25241.
981.0000000000,5547.0,2480.8,2688.1,25241.
982.0000000000,5547.0,2480.8,2688.2,25242.
983.0000000000,5547.1,2480.8,2686.3,25242.
984.0000000000,5547.1,2480.8,2686.3,25242.
985.0000000000,5547.1,2480.8,2685.5,25242.
986.0000000000,5547.2,2480.8,2685.8,25242.
987.0000000000,5547.2,2480.9,2686.4,25242.
988.0000000000,5547.2,2480.9,2686.9,25242.
989.0000000000,5547.3,2480.9,2687.4,25242.
990.0000000000,5547.3,2480.9,2687.8,25242.
991.0000000000,5547.3,2480.9,2688.2,25242.
992.0000000000,5547.4,2480.9,2688.5,25242.
993.0000000000,5547.4,2480.9,2688.8,25243.
994.0000000000,5547.4,2480.9,2689.0,25243.
995.0000000000,5547.5,2480.9,2689.2,25243.
996.0000000000,5547.5,2480.9,2689.4,25243.
997.0000000000,5547.5,2480.9,2689.6,25243.
998.0000000000,5547.6,2480.9,2689.7,25243.
999.0000000000,5547.6,2480.9,2689.8,25243.
1000.000000000,5547.6,2480.9,2689.1,25243.
1001.000000000,5547.7,2480.9,2689.2,25243.
1002.000000000,5547.7,2480.9,2689.4,25243.
1003.000000000,5547.7,2480.9,2689.6,25243.
1004.000000000,5547.8,2480.9,2689.8,25244.
1005.000000000,5547.8,2480.9,2690.0,25244.
1006.000000000,5547.8,2480.9,2690.2,25244.
1007.000000000,5547.9,2481.0,2690.4,25244.
1008.000000000,5547.9,2481.0,2690.6,25244.
1009.000000000,5547.9,2481.0,2690.7,25244.
1010.000000000,5548.0,2481.0,2690.8,25244.
1011.000000000,5548.0,2481.0,2690.9,25244.
1012.000000000,5548.0,2481.0,2681.3,25244.
1013.000000000,5548.1,2481.0,2679.3,25244.
1014.000000000,5548.1,2481.0,2680.4,25244.
1015.000000000,5548.1,2481.0,2682.1,25244.
1016.000000000,5548.2,2481.0,2683.8,25245.
1017.000000000,5548.2,2481.0,2685.3,25245.
1018.000000000,5548.2,2481.0,2686.6,25245.
1019.000000000,5548.3,2481.0,2687.6,25245.
1020.000000000,5548.3,2481.0,2688.5,25245.
1021.000000000,5548.3,2481.0,2689.2,25245.
1022.000000000,5548.4,2481.1,2689.8,25245.
1023.000000000,5548.4,2481.1,2690.3,25245.
1024.000000000,5548.4,2481.1,2690.7,25245.
1025.000000000,5548.5,2481.1,2690.4,25245.
1026.000000000,5548.5,2481.1,2689.6,25245.
1027.000000000,5548.5,2481.1,2669.6,25246.
1028.000000000,5548.6,2481.1,2660.1,25246.
1029.000000000,5548.6,2481.1,2662.2,25246.
1030.000000000,5548.6,2481.1,2666.4,25246.
1031.000000000,5548.7,2481.1,2670.9,25246.
1032.000000000,5548.7,2481.1,2674.9,25246.
1033.000000000,5548.7,2481.1,2677.5,25246.
1034.000000000,5548.8,2481.1,2668.5,25246.
1035.000000000,5548.8,2481.2,2670.2,25246.
1036.000000000,5548.8,2481.2,2673.4,25246.
1037.000000000,5548.9,2481.2,2676.7,25246.
1038.000000000,5548.9,2481.2,2679.7,25247.
1039.000000000,5549.0,2481.2,2682.1,25247.
1040.000000000,5549.0,2481.2,2684.2,25247.
1041.000000000,5549.0,2481.2,2685.4,25247.
1042.000000000,5549.1,2481.2,2686.2,25247.
1043.000000000,5549.1,2481.2,2687.3,25247.
1044.000000000,5549.1,2481.2,2688.3,25247.
1045.000000000,5549.2,2481.2,2689.2,25247.
1046.000000000,5549.2,2481.2,2689.9,25247.
1047.000000000,5549.2,2481.2,2690.5,25247.
1048.000000000,5549.3,2481.3,2690.7,25247.
1049.000000000,5549.3,2481.3,2690.3,25248.
1050.000000000,5549.3,2481.3,2690.4,25248.
1051.000000000,5549.4,2481.3,2690.6,25248.
1052.000000000,5549.4,2481.3,2691.0,25248.
1053.000000000,5549.4,2481.3,2691.4,25248.
1054.000000000,5549.5,2481.3,2691.8,25248.
1055.000000000,5549.5,2481.3,2692.1,25248.
1056.000000000,5549.5,2481.3,2692.4,25248.
1057.000000000,5549.6,2481.3,2692.6,25248.
1058.000000000,5549.6,2481.3,2692.9,25248.
1059.000000000,5549.6,2481.3,2693.1,25248.
1060.000000000,5549.7,2481.4,2692.9,25248.
1061.000000000,5549.7,2481.4,2691.2,25249.
1062.000000000,5549.8,2481.4,2684.0,25249.
1063.000000000,5549.8,2481.4,2683.6,25249.
1064.000000000,5549.8,2481.4,2684.8,25249.
1065.000000000,5549.9,2481.4,2686.3,25249.
1066.000000000,5549.9,2481.4,2687.8,25249.
1067.000000000,5549.9,2481.4,2689.0,25249.
1068.000000000,5550.0,2481.4,2690.1,25249.
1069.000000000,5550.0,2481.4,2691.0,25249.
1070.000000000,5550.0,2481.4,2691.7,25249.
1071.000000000,5550.1,2481.5,2692.3,25249.
1072.000000000,5550.1,2481.5,2692.8,25250.
1073.000000000,5550.1,2481.5,2693.2,25250.
1074.000000000,5550.2,2481.5,2693.5,25250.
1075.000000000,5550.2,2481.5,2693.8,25250.
1076.000000000,5550.2,2481.5,2694.1,25250.
1077.000000000,5550.3,2481.5,2685.7,25250.
1078.000000000,5550.3,2481.5,2685.4,25250.
1079.000000000,5550.4,2481.5,2686.5,25250.
1080.000000000,5550.4,2481.5,2687.9,25250.
1081.000000000,5550.4,2481.6,2689.2,25250.
1082.000000000,5550.5,2481.6,2690.4,25250.
1083.000000000,5550.5,2481.6,2691.4,25251.
1084.000000000,5550.5,2481.6,2692.2,25251.
1085.000000000,5550.6,2481.6,2692.9,25251.
1086.000000000,5550.6,2481.6,2693.5,25251.
1087.000000000,5550.6,2481.6,2694.0,25251.
1088.000000000,5550.7,2481.6,2694.4,25251.
1089.000000000,5550.7,2481.6,2694.7,25251.
1090.000000000,5550.8,2481.6,2695.0,25251.
1091.000000000,5550.8,2481.6,2687.9,25251.
1092.000000000,5550.8,2481.7,2686.2,25251.
1093.000000000,5550.9,2481.7,2687.1,25251.
1094.000000000,5550.9,2481.7,2688.5,25252.
1095.000000000,5550.9,2481.7,2689.8,25252.
1096.000000000,5551.0,2481.7,2691.1,25252.
1097.000000000,5551.0,2481.7,2692.0,25252.
1098.000000000,5551.1,2481.7,2691.6,25252.
1099.000000000,5551.1,2481.7,2692.2,25252.
1100.000000000,5551.1,2481.7,2693.0,25252.
1101.000000000,5551.2,2481.7,2693.7,25252.
1102.000000000,5551.2,2481.8,2694.3,25252.
1103.000000000,5551.2,2481.8,2694.8,25252.
1104.000000000,5551.3,2481.8,2695.3,25252.
1105.000000000,5551.3,2481.8,2695.6,25253.
1106.000000000,5551.4,2481.8,2696.0,25253.
1107.000000000,5551.4,2481.8,2696.2,25253.
1108.000000000,5551.4,2481.8,2696.5,25253.
1109.000000000,5551.5,2481.8,2696.7,25253.
1110.000000000,5551.5,2481.8,2696.8,25253.
1111.000000000,5551.5,2481.8,2697.0,25253.
1112.000000000,5551.6,2481.9,2697.1,25253.
1113.000000000,5551.6,2481.9,2697.3,25253.
1114.000000000,5551.6,2481.9,2697.4,25253.
1115.000000000,5551.7,2481.9,2697.5,25253.
1116.000000000,5551.7,2481.9,2697.6,25253.
1117.000000000,5551.8,2481.9,2697.8,25254.
1118.000000000,5551.8,2481.9,2697.9,25254.
1119.000000000,5551.8,2481.9,2698.0,25254.
1120.000000000,5551.9,2481.9,2698.1,25254.
1121.000000000,5551.9,2481.9,2698.2,25254.
1122.000000000,5551.9,2482.0,2693.8,25254.
1123.000000000,5552.0,2482.0,2693.6,25254.
1124.000000000,5552.0,2482.0,2694.2,25254.
1125.000000000,5552.1,2482.0,2695.0,25254.
1126.000000000,5552.1,2482.0,2695.7,25254.
1127.000000000,5552.1,2482.0,2696.3,25254.
1128.000000000,5552.2,2482.0,2696.9,25255.
1129.000000000,5552.2,2482.0,2697.3,25255.
1130.000000000,5552.3,2482.0,2697.7,25255.
1131.000000000,5552.3,2482.0,2698.1,25255.
1132.000000000,5552.3,2482.1,2698.4,25255.
1133.000000000,5552.4,2482.1,2698.6,25255.
1134.000000000,5552.4,2482.1,2698.8,25255.
1135.000000000,5552.4,2482.1,2699.0,25255.
1136.000000000,5552.5,2482.1,2699.2,25255.
1137.000000000,5552.5,2482.1,2699.3,25255.
1138.000000000,5552.6,2482.1,2699.5,25255.
1139.000000000,5552.6,2482.1,2699.6,25256.
1140.000000000,5552.6,2482.1,2699.7,25256.
1141.000000000,5552.7,2482.2,2699.8,25256.
1142.000000000,5552.7,2482.2,2700.0,25256.
1143.000000000,5552.7,2482.2,2700.1,25256.
1144.000000000,5552.8,2482.2,2700.2,25256.
1145.000000000,5552.8,2482.2,2700.3,25256.
1146.000000000,5552.9,2482.2,2700.4,25256.
1147.000000000,5552.9,2482.2,2700.5,25256.
1148.000000000,5552.9,2482.2,2698.9,25256.
1149.000000000,5553.0,2482.2,2694.1,25256.
1150.000000000,5553.0,2482.3,2694.2,25257.
1151.000000000,5553.0,2482.3,2695.0,25257.
1152.000000000,5553.1,2482.3,2696.0,25257.
1153.000000000,5553.1,2482.3,2697.0,25257.
1154.000000000,5553.2,2482.3,2697.8,25257.
1155.000000000,5553.2,2482.3,2698.6,25257.
1156.000000000,5553.2,2482.3,2699.2,25257.
1157.000000000,5553.3,2482.3,2699.7,25257.
1158.000000000,5553.3,2482.3,2700.1,25257.
1159.000000000,5553.4,2482.4,2700.4,25257.
1160.000000000,5553.4,2482.4,2700.7,25257.
1161.000000000,5553.4,2482.4,2701.0,25258.
1162.000000000,5553.5,2482.4,2701.2,25258.
1163.000000000,5553.5,2482.4,2693.6,25258.
1164.000000000,5553.5,2482.4,2688.3,25258.
1165.000000000,5553.6,2482.4,2681.6,25258.
1166.000000000,5553.6,2482.4,2675.6,25258.
1167.000000000,5553.7,2482.4,2673.5,25258.
1168.000000000,5553.7,2482.5,2676.9,25258.
1169.000000000,5553.7,2482.5,2681.0,25258.
1170.000000000,5553.8,2482.5,2684.9,25258.
1171.000000000,5553.8,2482.5,2688.2,25258.
1172.000000000,5553.9,2482.5,2690.8,25259.
1173.000000000,5553.9,2482.5,2693.1,25259.
1174.000000000,5553.9,2482.5,2691.3,25259.
1175.000000000,5554.0,2482.5,2692.6,25259.
1176.000000000,5554.0,2482.5,2694.2,25259.
1177.000000000,5554.0,2482.6,2695.7,25259.
1178.000000000,5554.1,2482.6,2697.0,25259.
1179.000000000,5554.1,2482.6,2697.6,25259.
1180.000000000,5554.2,2482.6,2698.5,25259.
1181.000000000,5554.2,2482.6,2699.3,25259.
1182.000000000,5554.2,2482.6,2700.0,25259.
1183.000000000,5554.3,2482.6,2700.5,25260.
1184.000000000,5554.3,2482.6,2701.0,25260.
1185.000000000,5554.3,2482.6,2701.4,25260.
1186.000000000,5554.4,2482.7,2701.8,25260.
1187.000000000,5554.4,2482.7,2702.0,25260.
1188.000000000,5554.5,2482.7,2702.2,25260.
1189.000000000,5554.5,2482.7,2702.4,25260.
1190.000000000,5554.5,2482.7,2702.6,25260.
1191.000000000,5554.6,2482.7,2702.8,25260.
1192.000000000,5554.6,2482.7,2703.0,25260.
1193.000000000,5554.6,2482.7,2703.1,25260.
1194.000000000,5554.7,2482.8,2703.3,25261.
1195.000000000,5554.7,2482.8,2703.4,25261.
1196.000000000,5554.8,2482.8,2703.5,25261.
1197.000000000,5554.8,2482.8,2703.5,25261.
1198.000000000,5554.8,2482.8,2703.6,25261.
1199.000000000,5554.9,2482.8,2700.5,25261.
1200.000000000,5554.9,2482.8,2700.4,25261.
1201.000000000,5555.0,2482.8,2700.9,25261.
1202.000000000,5555.0,2482.8,2701.5,25261.
1203.000000000,5555.0,2482.9,2680.6,25261.
1204.000000000,5555.1,2482.9,2675.1,25262.
1205.000000000,5555.1,2482.9,2677.5,25262.
1206.000000000,5555.1,2482.9,2681.4,25262.
1207.000000000,5555.2,2482.9,2685.4,25262.
1208.000000000,5555.2,2482.9,2688.9,25262.
1209.000000000,5555.3,2482.9,2691.9,25262.
1210.000000000,5555.3,2482.9,2694.1,25262.
1211.000000000,5555.3,2482.9,2696.1,25262.
1212.000000000,5555.4,2483.0,2697.8,25262.
1213.000000000,5555.4,2483.0,2697.1,25262.
1214.000000000,5555.5,2483.0,2698.1,25262.
1215.000000000,5555.5,2483.0,2699.2,25263.
1216.000000000,5555.5,2483.0,2700.2,25263.
1217.000000000,5555.6,2483.0,2701.1,25263.
1218.000000000,5555.6,2483.0,2701.8,25263.
1219.000000000,5555.7,2483.0,2702.4,25263.
1220.000000000,5555.7,2483.0,2703.0,25263.
1221.000000000,5555.7,2483.1,2703.4,25263.
1222.000000000,5555.8,2483.1,2703.8,25263.
1223.000000000,5555.8,2483.1,2704.1,25263.
1224.000000000,5555.9,2483.1,2704.4,25263.
1225.000000000,5555.9,2483.1,2703.9,25263.
1226.000000000,5555.9,2483.1,2704.1,25264.
1227.000000000,5556.0,2483.1,2704.4,25264.
1228.000000000,5556.0,2483.1,2704.6,25264.
1229.000000000,5556.1,2483.2,2704.8,25264.
1230.000000000,5556.1,2483.2,2705.0,25264.
1231.000000000,5556.2,2483.2,2704.1,25264.
1232.000000000,5556.2,2483.2,2703.5,25264.
1233.000000000,5556.2,2483.2,2703.7,25264.
1234.000000000,5556.3,2483.2,2701.5,25264.
1235.000000000,5556.3,2483.2,2694.9,25264.
1236.000000000,5556.4,2483.2,2693.8,25264.
1237.000000000,5556.4,2483.2,2695.2,25265.
1238.000000000,5556.4,2483.3,2697.0,25265.
1239.000000000,5556.5,2483.3,2698.7,25265.
1240.000000000,5556.5,2483.3,2700.2,25265.
1241.000000000,5556.6,2483.3,2701.5,25265.
1242.000000000,5556.6,2483.3,2702.6,25265.
1243.000000000,5556.6,2483.3,2703.4,25265.
1244.000000000,5556.7,2483.3,2704.1,25265.
1245.000000000,5556.7,2483.3,2704.7,25265.
1246.000000000,5556.8,2483.3,2704.8,25265.
1247.000000000,5556.8,2483.4,2705.2,25265.
1248.000000000,5556.8,2483.4,2704.8,25266.
1249.000000000,5556.9,2483.4,2691.1,25266.
1250.000000000,5556.9,2483.4,2687.6,25266.
1251.000000000,5557.0,2483.4,2689.1,25266.
1252.000000000,5557.0,2483.4,2691.7,25266.
1253.000000000,5557.0,2483.4,2694.4,25266.
1254.000000000,5557.1,2483.4,2696.9,25266.
1255.000000000,5557.1,2483.4,2698.9,25266.
1256.000000000,5557.2,2483.5,2700.6,25266.
1257.000000000,5557.2,2483.5,2702.0,25266.
1258.000000000,5557.2,2483.5,2703.2,25266.
1259.000000000,5557.3,2483.5,2704.1,25267.
1260.000000000,5557.3,2483.5,2704.7,25267.
1261.000000000,5557.4,2483.5,2705.3,25267.
1262.000000000,5557.4,2483.5,2705.8,25267.
1263.000000000,5557.4,2483.5,2706.2,25267.
1264.000000000,5557.5,2483.5,2706.6,25267.
1265.000000000,5557.5,2483.6,2706.9,25267.
1266.000000000,5557.6,2483.6,2707.2,25267.
1267.000000000,5557.6,2483.6,2704.3,25267.
1268.000000000,5557.6,2483.6,2704.3,25267.
1269.000000000,5557.7,2483.6,2704.8,25267.
1270.000000000,5557.7,2483.6,2705.5,25268.
1271.000000000,5557.8,2483.6,2706.0,25268.
1272.000000000,5557.8,2483.6,2706.6,25268.
1273.000000000,5557.8,2483.6,2704.0,25268.
1274.000000000,5557.9,2483.7,2680.9,25268.
1275.000000000,5557.9,2483.7,2679.4,25268.
1276.000000000,5558.0,2483.7,2682.3,25268.
1277.000000000,5558.0,2483.7,2686.4,25268.
1278.000000000,5558.0,2483.7,2690.4,25268.
1279.000000000,5558.1,2483.7,2693.9,25268.
1280.000000000,5558.1,2483.7,2696.8,25269.
1281.000000000,5558.2,2483.7,2699.2,25269.
1282.000000000,5558.2,2483.7,2701.2,25269.
1283.000000000,5558.3,2483.8,2702.7,25269.
1284.000000000,5558.3,2483.8,2704.0,25269.
1285.000000000,5558.3,2483.8,2705.0,25269.
1286.000000000,5558.4,2483.8,2705.9,25269.
1287.000000000,5558.4,2483.8,2706.5,25269.
1288.000000000,5558.5,2483.8,2707.1,25269.
1289.000000000,5558.5,2483.8,2707.5,25269.
1290.000000000,5558.5,2483.8,2707.9,25269.
1291.000000000,5558.6,2483.8,2708.2,25270.
1292.000000000,5558.6,2483.8,2708.5,25270.
1293.000000000,5558.7,2483.8,2708.8,25270.
1294.000000000,5558.7,2483.8,2709.0,25270.
1295.000000000,5558.7,2483.9,2709.1,25270.
1296.000000000,5558.8,2483.9,2709.3,25270.
1297.000000000,5558.8,2483.9,2709.5,25270.
1298.000000000,5558.9,2483.9,2709.6,25270.
1299.000000000,5558.9,2483.9,2709.7,25270.
1300.000000000,5558.9,2483.9,2709.8,25270.
1301.000000000,5559.0,2483.9,2710.0,25270.
1302.000000000,5559.0,2483.9,2710.1,25271.
1303.000000000,5559.1,2483.9,2710.1,25271.
1304.000000000,5559.1,2483.9,2707.7,25271.
1305.000000000,5559.1,2483.9,2707.5,25271.
1306.000000000,5559.2,2483.9,2707.8,25271.
1307.000000000,5559.2,2483.9,2708.2,25271.
1308.000000000,5559.3,2483.9,2708.7,25271.
1309.000000000,5559.3,2484.0,2709.1,25271.
1310.000000000,5559.3,2484.0,2709.5,25271.
1311.000000000,5559.4,2484.0,2709.9,25271.
1312.000000000,5559.4,2484.0,2710.2,25272.
1313.000000000,5559.5,2484.0,2710.4,25272.
1314.000000000,5559.5,2484.0,2710.6,25272.
1315.000000000,5559.5,2484.0,2710.8,25272.
1316.000000000,5559.6,2484.0,2711.0,25272.
1317.000000000,5559.6,2484.0,2711.2,25272.
1318.000000000,5559.7,2484.0,2711.3,25272.
1319.000000000,5559.7,2484.0,2711.5,25272.
1320.000000000,5559.7,2484.0,2711.6,25272.
1321.000000000,5559.8,2484.0,2703.1,25272.
1322.000000000,5559.8,2484.0,2695.3,25272.
1323.000000000,5559.9,2484.0,2693.1,25273.
1324.000000000,5559.9,2484.0,2694.5,25273.
1325.000000000,5559.9,2484.1,2691.9,25273.
1326.000000000,5560.0,2484.1,2692.7,25273.
1327.000000000,5560.0,2484.1,2694.9,25273.
1328.000000000,5560.0,2484.1,2679.8,25273.
1329.000000000,5560.1,2484.1,2679.2,25273.
1330.000000000,5560.1,2484.1,2679.8,25273.
1331.000000000,5560.2,2484.1,2680.1,25273.
1332.000000000,5560.2,2484.1,2684.6,25273.
1333.000000000,5560.2,2484.1,2688.8,25273.
1334.000000000,5560.3,2484.1,2693.0,25274.
1335.000000000,5560.3,2484.1,2696.6,25274.
1336.000000000,5560.4,2484.1,2699.4,25274.
1337.000000000,5560.4,2484.1,2700.5,25274.
1338.000000000,5560.4,2484.1,2701.9,25274.
1339.000000000,5560.5,2484.1,2702.4,25274.
1340.000000000,5560.5,2484.1,2703.2,25274.
1341.000000000,5560.6,2484.2,2703.9,25274.
1342.000000000,5560.6,2484.2,2702.6,25274.
1343.000000000,5560.6,2484.2,2703.7,25274.
1344.000000000,5560.7,2484.2,2705.1,25274.
1345.000000000,5560.7,2484.2,2706.4,25275.
1346.000000000,5560.8,2484.2,2707.5,25275.
1347.000000000,5560.8,2484.2,2708.5,25275.
1348.000000000,5560.8,2484.2,2709.3,25275.
1349.000000000,5560.9,2484.2,2709.9,25275.
1350.000000000,5560.9,2484.2,2709.6,25275.
1351.000000000,5561.0,2484.2,2710.0,25275.
1352.000000000,5561.0,2484.2,2708.1,25275.
1353.000000000,5561.0,2484.2,2708.2,25275.
1354.000000000,5561.1,2484.2,2707.7,25275.
1355.000000000,5561.1,2484.2,2708.4,25276.
1356.000000000,5561.2,2484.2,2709.2,25276.
1357.000000000,5561.2,2484.3,2709.9,25276.
1358.000000000,5561.2,2484.3,2710.5,25276.
1359.000000000,5561.3,2484.3,2711.1,25276.
1360.000000000,5561.3,2484.3,2711.5,25276.
1361.000000000,5561.4,2484.3,2711.9,25276.
1362.000000000,5561.4,2484.3,2712.2,25276.
1363.000000000,5561.4,2484.3,2712.5,25276.
1364.000000000,5561.5,2484.3,2701.4,25276.
1365.000000000,5561.5,2484.3,2675.2,25276.
1366.000000000,5561.6,2484.3,2672.2,25277.
1367.000000000,5561.6,2484.3,2676.6,25277.
1368.000000000,5561.6,2484.3,2682.4,25277.
1369.000000000,5561.7,2484.3,2688.0,25277.
1370.000000000,5561.7,2484.4,2692.8,25277.
1371.000000000,5561.8,2484.4,2696.9,25277.
1372.000000000,5561.8,2484.4,2700.2,25277.
1373.000000000,5561.8,2484.4,2702.9,25277.
1374.000000000,5561.9,2484.4,2705.0,25277.
1375.000000000,5561.9,2484.4,2706.7,25277.
1376.000000000,5562.0,2484.4,2708.1,25277.
1377.000000000,5562.0,2484.4,2709.2,25278.
1378.000000000,5562.0,2484.4,2710.1,25278.
1379.000000000,5562.1,2484.4,2710.8,25278.
1380.000000000,5562.1,2484.4,2711.4,25278.
1381.000000000,5562.2,2484.4,2711.9,25278.
1382.000000000,5562.2,2484.5,2712.3,25278.
1383.000000000,5562.2,2484.5,2712.7,25278.
1384.000000000,5562.3,2484.5,2713.0,25278.
1385.000000000,5562.3,2484.5,2713.2,25278.
1386.000000000,5562.4,2484.5,2713.4,25278.
1387.000000000,5562.4,2484.5,2713.6,25278.
1388.000000000,5562.4,2484.5,2713.8,25279.
1389.000000000,5562.5,2484.5,2713.9,25279.
1390.000000000,5562.5,2484.5,2714.0,25279.
1391.000000000,5562.6,2484.5,2714.1,25279.
1392.000000000,5562.6,2484.5,2714.3,25279.
1393.000000000,5562.7,2484.5,2714.4,25279.
1394.000000000,5562.7,2484.5,2714.5,25279.
1395.000000000,5562.7,2484.6,2714.6,25279.
1396.000000000,5562.8,2484.6,2714.7,25279.
1397.000000000,5562.8,2484.6,2714.8,25279.
1398.000000000,5562.9,2484.6,2714.9,25279.
1399.000000000,5562.9,2484.6,2715.0,25280.
1400.000000000,5562.9,2484.6,2715.1,25280.
1401.000000000,5563.0,2484.6,2715.2,25280.
1402.000000000,5563.0,2484.6,2715.3,25280.
1403.000000000,5563.1,2484.6,2715.4,25280.
1404.000000000,5563.1,2484.6,2710.5,25280.
1405.000000000,5563.1,2484.6,2710.1,25280.
1406.000000000,5563.2,2484.6,2710.7,25280.
1407.000000000,5563.2,2484.6,2710.8,25280.
1408.000000000,5563.3,2484.6,2711.6,25280.
1409.000000000,5563.3,2484.6,2712.4,25281.
1410.000000000,5563.3,2484.7,2705.7,25281.
1411.000000000,5563.4,2484.7,2705.7,25281.
1412.000000000,5563.4,2484.7,2707.0,25281.
1413.000000000,5563.5,2484.7,2708.5,25281.
1414.000000000,5563.5,2484.7,2710.0,25281.
1415.000000000,5563.6,2484.7,2711.2,25281.
1416.000000000,5563.6,2484.7,2712.3,25281.
1417.000000000,5563.6,2484.7,2713.2,25281.
1418.000000000,5563.7,2484.7,2713.9,25281.
1419.000000000,5563.7,2484.7,2714.5,25282.
1420.000000000,5563.8,2484.7,2715.0,25282.
1421.000000000,5563.8,2484.7,2715.4,25282.
1422.000000000,5563.8,2484.7,2715.7,25282.
1423.000000000,5563.9,2484.7,2716.0,25282.
1424.000000000,5563.9,2484.7,2716.3,25282.
1425.000000000,5564.0,2484.7,2716.5,25282.
1426.000000000,5564.0,2484.8,2716.0,25282.
1427.000000000,5564.0,2484.8,2716.1,25282.
1428.000000000,5564.1,2484.8,2716.3,25282.
1429.000000000,5564.1,2484.8,2716.6,25282.
1430.000000000,5564.2,2484.8,2716.8,25283.
1431.000000000,5564.2,2484.8,2717.0,25283.
1432.000000000,5564.2,2484.8,2717.2,25283.
1433.000000000,5564.3,2484.8,2714.5,25283.
1434.000000000,5564.3,2484.8,2709.7,25283.
1435.000000000,5564.4,2484.8,2693.6,25283.
1436.000000000,5564.4,2484.8,2692.2,25283.
1437.000000000,5564.4,2484.8,2695.0,25283.
1438.000000000,5564.5,2484.8,2698.7,25283.
1439.000000000,5564.5,2484.8,2702.2,25283.
1440.000000000,5564.6,2484.8,2705.2,25284.
1441.000000000,5564.6,2484.8,2707.8,25284.
1442.000000000,5564.6,2484.8,2709.9,25284.
1443.000000000,5564.7,2484.8,2711.2,25284.
1444.000000000,5564.7,2484.8,2712.5,25284.
1445.000000000,5564.8,2484.9,2713.7,25284.
1446.000000000,5564.8,2484.9,2714.5,25284.
1447.000000000,5564.8,2484.9,2715.3,25284.
1448.000000000,5564.9,2484.9,2715.9,25284.
1449.000000000,5564.9,2484.9,2716.5,25284.
1450.000000000,5565.0,2484.9,2716.9,25284.
1451.000000000,5565.0,2484.9,2717.3,25285.
1452.000000000,5565.0,2484.9,2717.2,25285.
1453.000000000,5565.1,2484.9,2717.5,25285.
1454.000000000,5565.1,2484.9,2717.1,25285.
1455.000000000,5565.1,2484.9,2717.3,25285.
1456.000000000,5565.2,2484.9,2717.6,25285.
1457.000000000,5565.2,2484.9,2717.9,25285.
1458.000000000,5565.3,2484.9,2718.2,25285.
1459.000000000,5565.3,2484.9,2718.4,25285.
1460.000000000,5565.3,2484.9,2718.5,25285.
1461.000000000,5565.4,2484.9,2718.6,25286.
1462.000000000,5565.4,2484.9,2718.8,25286.
1463.000000000,5565.5,2484.9,2718.6,25286.
1464.000000000,5565.5,2484.9,2718.7,25286.
1465.000000000,5565.5,2484.9,2718.9,25286.
1466.000000000,5565.6,2484.9,2719.1,25286.
1467.000000000,5565.6,2484.9,2719.3,25286.
1468.000000000,5565.6,2484.9,2719.5,25286.
1469.000000000,5565.7,2484.9,2719.6,25286.
1470.000000000,5565.7,2484.9,2719.8,25286.
1471.000000000,5565.8,2484.9,2719.9,25286.
1472.000000000,5565.8,2484.9,2720.0,25287.
1473.000000000,5565.8,2484.9,2720.2,25287.
1474.000000000,5565.9,2484.9,2720.3,25287.
1475.000000000,5565.9,2485.0,2719.8,25287.
1476.000000000,5565.9,2485.0,2718.6,25287.
1477.000000000,5566.0,2485.0,2716.0,25287.
1478.000000000,5566.0,2485.0,2716.2,25287.
1479.000000000,5566.1,2485.0,2713.4,25287.
1480.000000000,5566.1,2485.0,2713.9,25287.
1481.000000000,5566.1,2485.0,2715.0,25287.
1482.000000000,5566.2,2485.0,2716.1,25288.
1483.000000000,5566.2,2485.0,2717.0,25288.
1484.000000000,5566.2,2485.0,2717.9,25288.
1485.000000000,5566.3,2485.0,2718.6,25288.
1486.000000000,5566.3,2485.0,2719.2,25288.
1487.000000000,5566.4,2485.0,2719.7,25288.
1488.000000000,5566.4,2485.0,2720.1,25288.
1489.000000000,5566.4,2485.0,2720.3,25288.
1490.000000000,5566.5,2485.0,2720.5,25288.
1491.000000000,5566.5,2485.0,2720.8,25288.
1492.000000000,5566.5,2485.0,2721.0,25288.
1493.000000000,5566.6,2485.0,2721.3,25289.
1494.000000000,5566.6,2485.0,2721.4,25289.
1495.000000000,5566.7,2485.0,2721.6,25289.
1496.000000000,5566.7,2485.0,2721.8,25289.
1497.000000000,5566.7,2485.0,2721.8,25289.
1498.000000000,5566.8,2485.0,2721.9,25289.
1499.000000000,5566.8,2485.0,2722.1,25289.
1500.000000000,5566.8,2485.0,2722.2,25289.
1501.000000000,5566.9,2485.0,2722.3,25289.
1502.000000000,5566.9,2485.0,2722.4,25289.
1503.000000000,5567.0,2485.0,2722.6,25290.
1504.000000000,5567.0,2485.0,2722.7,25290.
1505.000000000,5567.0,2485.0,2722.8,25290.
1506.000000000,5567.1,2485.0,2711.8,25290.
1507.000000000,5567.1,2485.0,2711.3,25290.
1508.000000000,5567.1,2485.0,2712.6,25290.
1509.000000000,5567.2,2485.0,2714.1,25290.
1510.000000000,5567.2,2485.0,2715.7,25290.
1511.000000000,5567.3,2485.0,2717.2,25290.
1512.000000000,5567.3,2485.0,2717.0,25290.
1513.000000000,5567.3,2485.0,2717.9,25291.
1514.000000000,5567.4,2485.0,2718.9,25291.
1515.000000000,5567.4,2485.0,2719.9,25291.
1516.000000000,5567.4,2485.0,2720.6,25291.
1517.000000000,5567.5,2485.0,2721.3,25291.
1518.000000000,5567.5,2485.0,2721.8,25291.
1519.000000000,5567.6,2485.0,2722.3,25291.
1520.000000000,5567.6,2485.0,2722.7,25291.
1521.000000000,5567.6,2485.0,2723.0,25291.
1522.000000000,5567.7,2485.0,2723.3,25291.
1523.000000000,5567.7,2485.0,2723.5,25291.
1524.000000000,5567.7,2485.0,2723.7,25292.
1525.000000000,5567.8,2485.0,2723.1,25292.
1526.000000000,5567.8,2485.0,2723.3,25292.
1527.000000000,5567.9,2485.1,2723.5,25292.
1528.000000000,5567.9,2485.1,2723.7,25292.
1529.000000000,5567.9,2485.1,2724.0,25292.
1530.000000000,5568.0,2485.1,2724.2,25292.
1531.000000000,5568.0,2485.1,2724.2,25292.
1532.000000000,5568.0,2485.1,2724.3,25292.
1533.000000000,5568.1,2485.1,2724.5,25292.
1534.000000000,5568.1,2485.1,2724.7,25292.
1535.000000000,5568.2,2485.1,2724.8,25293.
1536.000000000,5568.2,2485.1,2725.0,25293.
1537.000000000,5568.2,2485.1,2725.1,25293.
1538.000000000,5568.3,2485.1,2725.2,25293.
1539.000000000,5568.3,2485.1,2725.4,25293.
1540.000000000,5568.3,2485.1,2725.5,25293.
1541.000000000,5568.4,2485.1,2725.6,25293.
1542.000000000,5568.4,2485.1,2725.7,25293.
1543.000000000,5568.5,2485.1,2725.8,25293.
1544.000000000,5568.5,2485.1,2725.8,25293.
1545.000000000,5568.5,2485.1,2725.9,25294.
1546.000000000,5568.6,2485.1,2726.0,25294.
1547.000000000,5568.6,2485.2,2726.1,25294.
1548.000000000,5568.6,2485.2,2726.2,25294.
1549.000000000,5568.7,2485.2,2721.4,25294.
1550.000000000,5568.7,2485.2,2721.3,25294.
1551.000000000,5568.8,2485.2,2721.9,25294.
1552.000000000,5568.8,2485.2,2722.7,25294.
1553.000000000,5568.8,2485.2,2714.2,25294.
1554.000000000,5568.9,2485.2,2714.4,25294.
1555.000000000,5568.9,2485.2,2716.0,25294.
1556.000000000,5568.9,2485.2,2717.8,25295.
1557.000000000,5569.0,2485.2,2719.5,25295.
1558.000000000,5569.0,2485.2,2721.0,25295.
1559.000000000,5569.1,2485.2,2722.3,25295.
1560.000000000,5569.1,2485.2,2723.3,25295.
1561.000000000,5569.1,2485.2,2724.2,25295.
1562.000000000,5569.2,2485.2,2721.8,25295.
1563.000000000,5569.2,2485.2,2721.4,25295.
1564.000000000,5569.2,2485.2,2721.1,25295.
1565.000000000,5569.3,2485.2,2717.8,25295.
1566.000000000,5569.3,2485.3,2718.6,25296.
1567.000000000,5569.4,2485.3,2719.6,25296.
1568.000000000,5569.4,2485.3,2719.6,25296.
1569.000000000,5569.4,2485.3,2720.8,25296.
1570.000000000,5569.5,2485.3,2722.1,25296.
1571.000000000,5569.5,2485.3,2723.2,25296.
1572.000000000,5569.5,2485.3,2724.2,25296.
1573.000000000,5569.6,2485.3,2725.0,25296.
1574.000000000,5569.6,2485.3,2725.7,25296.
1575.000000000,5569.7,2485.3,2726.2,25296.
1576.000000000,5569.7,2485.3,2726.7,25296.
1577.000000000,5569.7,2485.3,2727.1,25297.
1578.000000000,5569.8,2485.3,2727.4,25297.
1579.000000000,5569.8,2485.3,2727.7,25297.
1580.000000000,5569.8,2485.3,2727.9,25297.
1581.000000000,5569.9,2485.3,2728.1,25297.
1582.000000000,5569.9,2485.3,2728.3,25297.
1583.000000000,5570.0,2485.3,2728.5,25297.
1584.000000000,5570.0,2485.3,2728.6,25297.
1585.000000000,5570.0,2485.3,2728.7,25297.
1586.000000000,5570.1,2485.4,2728.9,25297.
1587.000000000,5570.1,2485.4,2729.0,25297.
1588.000000000,5570.2,2485.4,2729.1,25298.
1589.000000000,5570.2,2485.4,2729.2,25298.
1590.000000000,5570.2,2485.4,2729.3,25298.
1591.000000000,5570.3,2485.4,2729.4,25298.
1592.000000000,5570.3,2485.4,2725.7,25298.
1593.000000000,5570.4,2485.4,2725.5,25298.
1594.000000000,5570.4,2485.4,2726.1,25298.
1595.000000000,5570.4,2485.4,2726.7,25298.
1596.000000000,5570.5,2485.4,2727.3,25298.
1597.000000000,5570.5,2485.4,2727.9,25298.
1598.000000000,5570.5,2485.4,2728.3,25299.
1599.000000000,5570.6,2485.4,2728.7,25299.
1600.000000000,5570.6,2485.4,2729.1,25299.
1601.000000000,5570.7,2485.4,2721.8,25299.
1602.000000000,5570.7,2485.4,2721.2,25299.
1603.000000000,5570.7,2485.4,2716.0,25299.
1604.000000000,5570.8,2485.4,2716.9,25299.
1605.000000000,5570.8,2485.4,2718.6,25299.
1606.000000000,5570.9,2485.4,2720.7,25299.
1607.000000000,5570.9,2485.4,2722.6,25299.
1608.000000000,5570.9,2485.5,2724.2,25299.
1609.000000000,5571.0,2485.5,2725.6,25300.
1610.000000000,5571.0,2485.5,2719.1,25300.
1611.000000000,5571.1,2485.5,2719.4,25300.
1612.000000000,5571.1,2485.5,2696.3,25300.
1613.000000000,5571.1,2485.5,2693.7,25300.
1614.000000000,5571.2,2485.5,2697.2,25300.
1615.000000000,5571.2,2485.5,2700.7,25300.
1616.000000000,5571.2,2485.5,2701.4,25300.
1617.000000000,5571.3,2485.5,2705.2,25300.
1618.000000000,5571.3,2485.5,2709.6,25300.
1619.000000000,5571.4,2485.5,2713.6,25301.
1620.000000000,5571.4,2485.5,2716.9,25301.
1621.000000000,5571.4,2485.5,2719.7,25301.
1622.000000000,5571.5,2485.5,2722.0,25301.
1623.000000000,5571.5,2485.5,2723.8,25301.
1624.000000000,5571.6,2485.5,2725.2,25301.
1625.000000000,5571.6,2485.5,2726.4,25301.
1626.000000000,5571.6,2485.5,2727.4,25301.
1627.000000000,5571.7,2485.5,2728.1,25301.
1628.000000000,5571.7,2485.5,2728.7,25301.
1629.000000000,5571.7,2485.5,2729.2,25301.
1630.000000000,5571.8,2485.5,2729.7,25301.
1631.000000000,5571.8,2485.5,2730.0,25302.
1632.000000000,5571.8,2485.5,2730.3,25302.
1633.000000000,5571.9,2485.5,2730.6,25302.
1634.000000000,5571.9,2485.5,2730.8,25302.
1635.000000000,5572.0,2485.5,2731.0,25302.
1636.000000000,5572.0,2485.5,2731.1,25302.
1637.000000000,5572.0,2485.5,2731.2,25302.
1638.000000000,5572.1,2485.5,2731.3,25302.
1639.000000000,5572.1,2485.5,2729.4,25302.
1640.000000000,5572.1,2485.5,2729.0,25302.
1641.000000000,5572.2,2485.5,2729.3,25303.
1642.000000000,5572.2,2485.5,2729.8,25303.
1643.000000000,5572.2,2485.5,2730.3,25303.
1644.000000000,5572.3,2485.5,2730.7,25303.
1645.000000000,5572.3,2485.5,2731.0,25303.
1646.000000000,5572.4,2485.5,2731.4,25303.
1647.000000000,5572.4,2485.5,2731.4,25303.
1648.000000000,5572.4,2485.5,2731.3,25303.
1649.000000000,5572.5,2485.5,2728.6,25303.
1650.000000000,5572.5,2485.5,2725.1,25303.
1651.000000000,5572.5,2485.5,2725.4,25303.
1652.000000000,5572.6,2485.5,2726.4,25304.
1653.000000000,5572.6,2485.5,2727.6,25304.
1654.000000000,5572.6,2485.5,2728.6,25304.
1655.000000000,5572.7,2485.5,2729.5,25304.
1656.000000000,5572.7,2485.5,2729.6,25304.
1657.000000000,5572.7,2485.5,2728.9,25304.
1658.000000000,5572.8,2485.6,2727.4,25304.
1659.000000000,5572.8,2485.6,2727.0,25304.
1660.000000000,5572.9,2485.6,2727.3,25304.
1661.000000000,5572.9,2485.6,2727.9,25304.
1662.000000000,5572.9,2485.6,2728.9,25304.
1663.000000000,5573.0,2485.6,2729.8,25305.
1664.000000000,5573.0,2485.6,2730.6,25305.
1665.000000000,5573.0,2485.6,2731.2,25305.
1666.000000000,5573.1,2485.6,2724.5,25305.
1667.000000000,5573.1,2485.6,2724.5,25305.
1668.000000000,5573.1,2485.6,2725.7,25305.
1669.000000000,5573.2,2485.6,2727.1,25305.
1670.000000000,5573.2,2485.6,2728.4,25305.
1671.000000000,5573.2,2485.6,2729.6,25305.
1672.000000000,5573.3,2485.6,2730.5,25305.
1673.000000000,5573.3,2485.6,2730.4,25306.
1674.000000000,5573.3,2485.6,2730.6,25306.
1675.000000000,5573.4,2485.6,2730.0,25306.
1676.000000000,5573.4,2485.6,2729.1,25306.
1677.000000000,5573.4,2485.6,2729.7,25306.
1678.000000000,5573.5,2485.6,2730.4,25306.
1679.000000000,5573.5,2485.6,2731.2,25306.
1680.000000000,5573.5,2485.6,2731.9,25306.
1681.000000000,5573.6,2485.6,2732.1,25306.
1682.000000000,5573.6,2485.6,2723.2,25306.
1683.000000000,5573.6,2485.6,2723.2,25306.
1684.000000000,5573.7,2485.6,2724.5,25307.
1685.000000000,5573.7,2485.6,2726.2,25307.
1686.000000000,5573.8,2485.6,2727.9,25307.
1687.000000000,5573.8,2485.6,2729.3,25307.
1688.000000000,5573.8,2485.6,2730.5,25307.
1689.000000000,5573.9,2485.6,2730.8,25307.
1690.000000000,5573.9,2485.6,2731.3,25307.
1691.000000000,5573.9,2485.6,2732.0,25307.
1692.000000000,5574.0,2485.6,2732.7,25307.
1693.000000000,5574.0,2485.6,2733.3,25307.
1694.000000000,5574.0,2485.6,2733.8,25307.
1695.000000000,5574.1,2485.6,2734.2,25307.
1696.000000000,5574.1,2485.6,2734.6,25308.
1697.000000000,5574.1,2485.6,2732.6,25308.
1698.000000000,5574.2,2485.6,2729.9,25308.
1699.000000000,5574.2,2485.6,2729.9,25308.
1700.000000000,5574.2,2485.6,2728.9,25308.
1701.000000000,5574.3,2485.6,2729.7,25308.
1702.000000000,5574.3,2485.6,2730.8,25308.
1703.000000000,5574.3,2485.6,2731.8,25308.
1704.000000000,5574.4,2485.6,2732.7,25308.
1705.000000000,5574.4,2485.6,2733.5,25308.
1706.000000000,5574.4,2485.6,2734.2,25308.
1707.000000000,5574.5,2485.6,2734.7,25309.
1708.000000000,5574.5,2485.6,2735.0,25309.
1709.000000000,5574.5,2485.6,2735.4,25309.
1710.000000000,5574.6,2485.6,2735.7,25309.
1711.000000000,5574.6,2485.6,2735.9,25309.
1712.000000000,5574.6,2485.6,2736.2,25309.
1713.000000000,5574.7,2485.6,2736.4,25309.
1714.000000000,5574.7,2485.6,2736.6,25309.
1715.000000000,5574.7,2485.6,2736.8,25309.
1716.000000000,5574.8,2485.6,2736.9,25309.
1717.000000000,5574.8,2485.6,2737.1,25309.
1718.000000000,5574.8,2485.6,2737.2,25310.
1719.000000000,5574.9,2485.6,2737.3,25310.
1720.000000000,5574.9,2485.6,2737.5,25310.
1721.000000000,5574.9,2485.6,2737.6,25310.
1722.000000000,5575.0,2485.6,2737.7,25310.
1723.000000000,5575.0,2485.7,2737.8,25310.
1724.000000000,5575.0,2485.7,2737.7,25310.
1725.000000000,5575.1,2485.7,2737.8,25310.
1726.000000000,5575.1,2485.7,2737.9,25310.
1727.000000000,5575.1,2485.7,2737.9,25310.
1728.000000000,5575.2,2485.7,2738.0,25310.
1729.000000000,5575.2,2485.7,2730.0,25311.
1730.000000000,5575.2,2485.7,2724.8,25311.
1731.000000000,5575.3,2485.7,2709.2,25311.
1732.000000000,5575.3,2485.7,2694.1,25311.
1733.000000000,5575.3,2485.7,2689.7,25311.
1734.000000000,5575.4,2485.7,2692.9,25311.
1735.000000000,5575.4,2485.7,2698.9,25311.
1736.000000000,5575.4,2485.7,2705.6,25311.
1737.000000000,5575.5,2485.7,2711.7,25311.
1738.000000000,5575.5,2485.7,2712.1,25311.
1739.000000000,5575.5,2485.7,2715.3,25311.
1740.000000000,5575.6,2485.7,2719.2,25312.
1741.000000000,5575.6,2485.7,2722.8,25312.
1742.000000000,5575.6,2485.7,2725.7,25312.
1743.000000000,5575.7,2485.7,2728.2,25312.
1744.000000000,5575.7,2485.7,2727.7,25312.
1745.000000000,5575.7,2485.7,2729.0,25312.
1746.000000000,5575.8,2485.7,2730.6,25312.
1747.000000000,5575.8,2485.7,2732.0,25312.
1748.000000000,5575.8,2485.7,2733.2,25312.
1749.000000000,5575.9,2485.7,2734.3,25312.
1750.000000000,5575.9,2485.7,2735.0,25312.
1751.000000000,5575.9,2485.7,2735.7,25312.
1752.000000000,5576.0,2485.7,2736.3,25313.
1753.000000000,5576.0,2485.7,2736.8,25313.
1754.000000000,5576.0,2485.7,2737.2,25313.
1755.000000000,5576.1,2485.7,2737.5,25313.
1756.000000000,5576.1,2485.7,2737.8,25313.
1757.000000000,5576.1,2485.7,2738.0,25313.
1758.000000000,5576.2,2485.7,2738.2,25313.
1759.000000000,5576.2,2485.7,2738.4,25313.
1760.000000000,5576.2,2485.7,2738.6,25313.
1761.000000000,5576.3,2485.7,2738.7,25313.
1762.000000000,5576.3,2485.7,2738.8,25313.
1763.000000000,5576.3,2485.7,2739.0,25314.
1764.000000000,5576.4,2485.7,2739.1,25314.
1765.000000000,5576.4,2485.7,2739.2,25314.
1766.000000000,5576.4,2485.7,2739.3,25314.
1767.000000000,5576.5,2485.7,2739.4,25314.
1768.000000000,5576.5,2485.7,2739.5,25314.
1769.000000000,5576.5,2485.7,2739.6,25314.
1770.000000000,5576.5,2485.7,2739.7,25314.
1771.000000000,5576.6,2485.7,2739.8,25314.
1772.000000000,5576.6,2485.7,2739.9,25314.
1773.000000000,5576.6,2485.7,2739.9,25314.
1774.000000000,5576.7,2485.7,2739.9,25314.
1775.000000000,5576.7,2485.7,2740.0,25315.
1776.000000000,5576.7,2485.7,2740.1,25315.
1777.000000000,5576.8,2485.7,2739.5,25315.
1778.000000000,5576.8,2485.7,2739.5,25315.
1779.000000000,5576.8,2485.7,2739.5,25315.
1780.000000000,5576.9,2485.7,2739.7,25315.
1781.000000000,5576.9,2485.7,2739.9,25315.
1782.000000000,5576.9,2485.7,2740.1,25315.
1783.000000000,5577.0,2485.7,2740.3,25315.
1784.000000000,5577.0,2485.7,2740.5,25315.
1785.000000000,5577.0,2485.7,2740.7,25315.
1786.000000000,5577.1,2485.7,2740.8,25316.
1787.000000000,5577.1,2485.7,2741.0,25316.
1788.000000000,5577.1,2485.7,2741.1,25316.
1789.000000000,5577.2,2485.7,2741.2,25316.
1790.000000000,5577.2,2485.7,2741.3,25316.
1791.000000000,5577.2,2485.7,2741.4,25316.
1792.000000000,5577.3,2485.7,2741.5,25316.
1793.000000000,5577.3,2485.7,2741.6,25316.
1794.000000000,5577.3,2485.7,2741.7,25316.
1795.000000000,5577.4,2485.7,2741.8,25316.
1796.000000000,5577.4,2485.7,2741.9,25316.
1797.000000000,5577.4,2485.7,2742.0,25316.
1798.000000000,5577.5,2485.7,2742.1,25317.
1799.000000000,5577.5,2485.7,2742.2,25317.
1800.000000000,5577.5,2485.7,2742.3,25317.
1801.000000000,5577.6,2485.7,2740.2,25317.
1802.000000000,5577.6,2485.7,2732.2,25317.
1803.000000000,5577.7,2485.7,2729.8,25317.
1804.000000000,5577.7,2485.7,2731.0,25317.
1805.000000000,5577.7,2485.7,2732.7,25317.
1806.000000000,5577.8,2485.7,2734.5,25317.
1807.000000000,5577.8,2485.7,2736.1,25317.
1808.000000000,5577.8,2485.7,2737.5,25317.
1809.000000000,5577.9,2485.7,2738.6,25318.
1810.000000000,5577.9,2485.7,2739.6,25318.
1811.000000000,5577.9,2485.7,2740.0,25318.
1812.000000000,5578.0,2485.7,2737.8,25318.
1813.000000000,5578.0,2485.7,2738.1,25318.
1814.000000000,5578.0,2485.7,2738.3,25318.
1815.000000000,5578.1,2485.7,2739.1,25318.
1816.000000000,5578.1,2485.7,2739.9,25318.
1817.000000000,5578.1,2485.7,2740.6,25318.
1818.000000000,5578.2,2485.7,2741.1,25318.
1819.000000000,5578.2,2485.7,2741.7,25318.
1820.000000000,5578.2,2485.7,2742.1,25319.
1821.000000000,5578.3,2485.7,2742.5,25319.
1822.000000000,5578.3,2485.7,2742.5,25319.
1823.000000000,5578.3,2485.7,2742.6,25319.
1824.000000000,5578.4,2485.7,2742.8,25319.
1825.000000000,5578.4,2485.7,2743.1,25319.
1826.000000000,5578.4,2485.7,2743.3,25319.
1827.000000000,5578.5,2485.7,2743.5,25319.
1828.000000000,5578.5,2485.7,2743.7,25319.
1829.000000000,5578.5,2485.7,2743.8,25319.
1830.000000000,5578.6,2485.7,2744.0,25319.
1831.000000000,5578.6,2485.7,2744.2,25319.
1832.000000000,5578.6,2485.7,2744.3,25320.
1833.000000000,5578.6,2485.7,2744.5,25320.
1834.000000000,5578.7,2485.7,2744.6,25320.
1835.000000000,5578.7,2485.7,2744.7,25320.
1836.000000000,5578.7,2485.7,2744.8,25320.
1837.000000000,5578.8,2485.7,2744.9,25320.
1838.000000000,5578.8,2485.7,2745.1,25320.
1839.000000000,5578.8,2485.7,2745.2,25320.
1840.000000000,5578.9,2485.7,2745.3,25320.
1841.000000000,5578.9,2485.7,2745.4,25320.
1842.000000000,5578.9,2485.7,2745.3,25320.
1843.000000000,5579.0,2485.7,2745.4,25320.
1844.000000000,5579.0,2485.8,2745.5,25321.
1845.000000000,5579.0,2485.8,2745.5,25321.
1846.000000000,5579.1,2485.8,2745.5,25321.
1847.000000000,5579.1,2485.8,2745.6,25321.
1848.000000000,5579.1,2485.8,2745.7,25321.
1849.000000000,5579.2,2485.8,2745.9,25321.
1850.000000000,5579.2,2485.8,2746.0,25321.
1851.000000000,5579.2,2485.8,2746.1,25321.
1852.000000000,5579.3,2485.8,2746.3,25321.
1853.000000000,5579.3,2485.8,2746.4,25321.
1854.000000000,5579.3,2485.8,2746.5,25321.
1855.000000000,5579.4,2485.8,2746.6,25321.
1856.000000000,5579.4,2485.8,2746.7,25322.
1857.000000000,5579.4,2485.8,2746.8,25322.
1858.000000000,5579.5,2485.8,2746.9,25322.
1859.000000000,5579.5,2485.8,2747.0,25322.
1860.000000000,5579.5,2485.8,2746.9,25322.
1861.000000000,5579.6,2485.8,2747.0,25322.
1862.000000000,5579.6,2485.8,2747.1,25322.
1863.000000000,5579.6,2485.8,2747.2,25322.
1864.000000000,5579.7,2485.8,2747.3,25322.
1865.000000000,5579.7,2485.8,2747.4,25322.
1866.000000000,5579.7,2485.8,2747.5,25322.
1867.000000000,5579.8,2485.8,2747.6,25322.
1868.000000000,5579.8,2485.8,2747.7,25323.
1869.000000000,5579.8,2485.8,2747.8,25323.
1870.000000000,5579.9,2485.8,2747.4,25323.
1871.000000000,5579.9,2485.8,2747.3,25323.
1872.000000000,5579.9,2485.8,2747.4,25323.
1873.000000000,5580.0,2485.8,2747.6,25323.
1874.000000000,5580.0,2485.8,2747.8,25323.
1875.000000000,5580.0,2485.9,2748.0,25323.
1876.000000000,5580.1,2485.9,2747.4,25323.
1877.000000000,5580.1,2485.9,2745.2,25323.
1878.000000000,5580.2,2485.9,2736.0,25323.
1879.000000000,5580.2,2485.9,2735.3,25324.
1880.000000000,5580.2,2485.9,2736.8,25324.
1881.000000000,5580.3,2485.9,2738.6,25324.
1882.000000000,5580.3,2485.9,2740.4,25324.
1883.000000000,5580.3,2485.9,2742.1,25324.
1884.000000000,5580.4,2485.9,2743.5,25324.
1885.000000000,5580.4,2485.9,2744.7,25324.
1886.000000000,5580.4,2485.9,2745.2,25324.
1887.000000000,5580.5,2485.9,2745.9,25324.
1888.000000000,5580.5,2485.9,2746.6,25324.
1889.000000000,5580.5,2485.9,2747.2,25324.
1890.000000000,5580.6,2485.9,2747.7,25324.
1891.000000000,5580.6,2485.9,2748.1,25324.
1892.000000000,5580.6,2485.9,2748.5,25325.
1893.000000000,5580.7,2486.0,2748.8,25325.
1894.000000000,5580.7,2486.0,2749.1,25325.
1895.000000000,5580.7,2486.0,2749.3,25325.
1896.000000000,5580.8,2486.0,2749.5,25325.
1897.000000000,5580.8,2486.0,2749.7,25325.
1898.000000000,5580.8,2486.0,2749.8,25325.
1899.000000000,5580.9,2486.0,2750.0,25325.
1900.000000000,5580.9,2486.0,2750.1,25325.
1901.000000000,5581.0,2486.0,2750.2,25325.
1902.000000000,5581.0,2486.0,2750.3,25325.
1903.000000000,5581.0,2486.0,2750.5,25325.
1904.000000000,5581.1,2486.0,2750.6,25326.
1905.000000000,5581.1,2486.0,2750.7,25326.
1906.000000000,5581.1,2486.0,2750.8,25326.
1907.000000000,5581.2,2486.0,2750.9,25326.
1908.000000000,5581.2,2486.0,2751.0,25326.
1909.000000000,5581.2,2486.0,2751.1,25326.
1910.000000000,5581.3,2486.0,2751.2,25326.
1911.000000000,5581.3,2486.0,2751.2,25326.
1912.000000000,5581.3,2486.0,2751.3,25326.
1913.000000000,5581.4,2486.0,2751.0,25326.
1914.000000000,5581.4,2486.1,2751.0,25326.
1915.000000000,5581.4,2486.1,2751.2,25326.
1916.000000000,5581.5,2486.1,2751.3,25327.
1917.000000000,5581.5,2486.1,2751.5,25327.
1918.000000000,5581.5,2486.1,2751.6,25327.
1919.000000000,5581.6,2486.1,2751.8,25327.
1920.000000000,5581.6,2486.1,2751.9,25327.
1921.000000000,5581.6,2486.1,2752.0,25327.
1922.000000000,5581.7,2486.1,2752.1,25327.
1923.000000000,5581.7,2486.1,2752.3,25327.
1924.000000000,5581.7,2486.1,2752.4,25327.
1925.000000000,5581.8,2486.1,2752.5,25327.
1926.000000000,5581.8,2486.1,2752.6,25327.
1927.000000000,5581.8,2486.1,2752.7,25327.
1928.000000000,5581.9,2486.1,2752.8,25328.
1929.000000000,5581.9,2486.1,2752.9,25328.
1930.000000000,5581.9,2486.1,2752.7,25328.
1931.000000000,5582.0,2486.1,2752.8,25328.
1932.000000000,5582.0,2486.1,2752.9,25328.
1933.000000000,5582.0,2486.1,2753.0,25328.
1934.000000000,5582.1,2486.1,2753.2,25328.
1935.000000000,5582.1,2486.1,2753.3,25328.
1936.000000000,5582.1,2486.2,2753.4,25328.
1937.000000000,5582.2,2486.2,2753.5,25328.
1938.000000000,5582.2,2486.2,2753.5,25328.
1939.000000000,5582.2,2486.2,2753.6,25328.
1940.000000000,5582.3,2486.2,2753.7,25329.
1941.000000000,5582.3,2486.2,2753.8,25329.
1942.000000000,5582.3,2486.2,2752.4,25329.
1943.000000000,5582.4,2486.2,2752.4,25329.
1944.000000000,5582.4,2486.2,2752.7,25329.
1945.000000000,5582.4,2486.2,2753.1,25329.
1946.000000000,5582.5,2486.2,2753.4,25329.
1947.000000000,5582.5,2486.2,2753.7,25329.
1948.000000000,5582.5,2486.2,2753.9,25329.
1949.000000000,5582.6,2486.2,2753.7,25329.
1950.000000000,5582.6,2486.2,2743.3,25329.
1951.000000000,5582.6,2486.2,2741.2,25329.
1952.000000000,5582.7,2486.2,2742.5,25330.
1953.000000000,5582.7,2486.2,2744.4,25330.
1954.000000000,5582.8,2486.2,2746.3,25330.
1955.000000000,5582.8,2486.2,2748.0,25330.
1956.000000000,5582.8,2486.2,2749.5,25330.
1957.000000000,5582.9,2486.2,2750.7,25330.
1958.000000000,5582.9,2486.2,2751.7,25330.
1959.000000000,5582.9,2486.2,2752.5,25330.
1960.000000000,5583.0,2486.3,2753.1,25330.
1961.000000000,5583.0,2486.3,2753.7,25330.
1962.000000000,5583.0,2486.3,2754.1,25330.
1963.000000000,5583.1,2486.3,2754.5,25330.
1964.000000000,5583.1,2486.3,2754.8,25331.
1965.000000000,5583.1,2486.3,2755.0,25331.
1966.000000000,5583.2,2486.3,2754.3,25331.
1967.000000000,5583.2,2486.3,2744.2,25331.
1968.000000000,5583.2,2486.3,2743.7,25331.
1969.000000000,5583.3,2486.3,2745.1,25331.
1970.000000000,5583.3,2486.3,2746.9,25331.
1971.000000000,5583.3,2486.3,2748.6,25331.
1972.000000000,5583.4,2486.3,2750.1,25331.
1973.000000000,5583.4,2486.3,2751.4,25331.
1974.000000000,5583.4,2486.3,2752.5,25331.
1975.000000000,5583.5,2486.3,2753.3,25331.
1976.000000000,5583.5,2486.3,2754.1,25332.
1977.000000000,5583.5,2486.3,2754.6,25332.
1978.000000000,5583.6,2486.3,2755.1,25332.
1979.000000000,5583.6,2486.3,2755.5,25332.
1980.000000000,5583.6,2486.3,2755.9,25332.
1981.000000000,5583.7,2486.3,2755.6,25332.
1982.000000000,5583.7,2486.3,2755.8,25332.
1983.000000000,5583.7,2486.3,2756.1,25332.
1984.000000000,5583.8,2486.3,2756.3,25332.
1985.000000000,5583.8,2486.3,2756.6,25332.
1986.000000000,5583.8,2486.4,2756.8,25332.
1987.000000000,5583.9,2486.4,2757.0,25332.
1988.000000000,5583.9,2486.4,2757.2,25333.
1989.000000000,5583.9,2486.4,2757.3,25333.
1990.000000000,5584.0,2486.4,2757.5,25333.
1991.000000000,5584.0,2486.4,2757.6,25333.
1992.000000000,5584.0,2486.4,2757.7,25333.
1993.000000000,5584.1,2486.4,2757.8,25333.
1994.000000000,5584.1,2486.4,2758.0,25333.
1995.000000000,5584.1,2486.4,2758.0,25333.
1996.000000000,5584.2,2486.4,2757.4,25333.
1997.000000000,5584.2,2486.4,2757.5,25333.
1998.000000000,5584.2,2486.4,2757.7,25333.
1999.000000000,5584.3,2486.4,2757.7,25333.
2000.000000000,5584.3,2486.4,2757.9,25334.
2001.000000000,5584.3,2486.4,2758.1,25334.
2002.000000000,5584.4,2486.4,2758.3,25334.
2003.000000000,5584.4,2486.4,2758.5,25334.
2004.000000000,5584.4,2486.4,2758.7,25334.
2005.000000000,5584.5,2486.4,2758.8,25334.
2006.000000000,5584.5,2486.4,2758.9,25334.
2007.000000000,5584.5,2486.4,2758.5,25334.
2008.000000000,5584.6,2486.4,2758.6,25334.
2009.000000000,5584.6,2486.5,2758.7,25334.
2010.000000000,5584.6,2486.5,2758.9,25334.
2011.000000000,5584.7,2486.5,2759.1,25334.
2012.000000000,5584.7,2486.5,2758.2,25335.
2013.000000000,5584.7,2486.5,2756.5,25335.
2014.000000000,5584.8,2486.5,2752.3,25335.
2015.000000000,5584.8,2486.5,2747.9,25335.
2016.000000000,5584.8,2486.5,2746.7,25335.
2017.000000000,5584.9,2486.5,2745.0,25335.
2018.000000000,5584.9,2486.5,2746.8,25335.
2019.000000000,5584.9,2486.5,2749.0,25335.
2020.000000000,5585.0,2486.5,2751.1,25335.
2021.000000000,5585.0,2486.5,2752.9,25335.
2022.000000000,5585.0,2486.5,2754.4,25335.
2023.000000000,5585.1,2486.5,2755.6,25335.
2024.000000000,5585.1,2486.5,2756.7,25335.
2025.000000000,5585.1,2486.5,2757.5,25336.
2026.000000000,5585.2,2486.5,2758.2,25336.
2027.000000000,5585.2,2486.5,2758.7,25336.
2028.000000000,5585.2,2486.5,2759.2,25336.
2029.000000000,5585.3,2486.5,2759.6,25336.
2030.000000000,5585.3,2486.6,2759.9,25336.
2031.000000000,5585.3,2486.6,2760.2,25336.
2032.000000000,5585.4,2486.6,2760.4,25336.
2033.000000000,5585.4,2486.6,2760.6,25336.
2034.000000000,5585.4,2486.6,2760.8,25336.
2035.000000000,5585.5,2486.6,2761.0,25336.
2036.000000000,5585.5,2486.6,2761.1,25336.
2037.000000000,5585.5,2486.6,2761.2,25336.
2038.000000000,5585.6,2486.6,2750.9,25337.
2039.000000000,5585.6,2486.6,2750.1,25337.
2040.000000000,5585.7,2486.6,2751.4,25337.
2041.000000000,5585.7,2486.6,2753.0,25337.
2042.000000000,5585.7,2486.6,2754.6,25337.
2043.000000000,5585.8,2486.6,2756.1,25337.
2044.000000000,5585.8,2486.6,2757.3,25337.
2045.000000000,5585.8,2486.6,2758.3,25337.
2046.000000000,5585.9,2486.6,2759.1,25337.
2047.000000000,5585.9,2486.6,2759.8,25337.
2048.000000000,5585.9,2486.6,2760.3,25337.
2049.000000000,5586.0,2486.6,2756.7,25337.
2050.000000000,5586.0,2486.6,2754.1,25338.
2051.000000000,5586.0,2486.6,2751.1,25338.
2052.000000000,5586.1,2486.6,2751.1,25338.
2053.000000000,5586.1,2486.7,2752.7,25338.
2054.000000000,5586.1,2486.7,2754.4,25338.
2055.000000000,5586.2,2486.7,2756.0,25338.
2056.000000000,5586.2,2486.7,2757.3,25338.
2057.000000000,5586.2,2486.7,2758.4,25338.
2058.000000000,5586.3,2486.7,2758.5,25338.
2059.000000000,5586.3,2486.7,2757.5,25338.
2060.000000000,5586.3,2486.7,2758.2,25338.
2061.000000000,5586.4,2486.7,2759.0,25338.
2062.000000000,5586.4,2486.7,2759.8,25339.
2063.000000000,5586.4,2486.7,2760.5,25339.
2064.000000000,5586.5,2486.7,2761.1,25339.
2065.000000000,5586.5,2486.7,2761.6,25339.
2066.000000000,5586.5,2486.7,2762.0,25339.
2067.000000000,5586.6,2486.7,2762.4,25339.
2068.000000000,5586.6,2486.7,2762.7,25339.
2069.000000000,5586.6,2486.7,2762.9,25339.
