time,FINEGAN,704,703,DOLAN,701
1.000000000000,-106.32,-12.776,-11.175,-15331.,-17887.
2.000000000000,-106.28,-12.774,-11.172,-15332.,-17891.
3.000000000000,-106.25,-12.775,-11.171,-15333.,-17893.
4.000000000000,-106.33,-12.791,-11.184,-15333.,-17896.
5.000000000000,-106.32,-12.797,-11.187,-15334.,-17899.
6.000000000000,-106.26,-12.796,-11.184,-15335.,-17902.
7.000000000000,-106.23,-12.797,-11.183,-15336.,-17905.
8.000000000000,-106.21,-12.799,-11.183,-15337.,-17908.
9.000000000000,-106.81,-12.874,-11.255,-15339.,-17912.
10.00000000000,-107.24,-12.935,-11.314,-15340.,-17916.
11.00000000000,-106.83,-12.894,-11.271,-15341.,-17920.
12.00000000000,-106.67,-12.871,-11.244,-15342.,-17923.
13.00000000000,-106.58,-12.857,-11.230,-15343.,-17926.
14.00000000000,-106.51,-12.850,-11.222,-15344.,-17928.
15.00000000000,-106.46,-12.847,-11.218,-15345.,-17931.
16.00000000000,-106.42,-12.845,-11.216,-15346.,-17933.
17.00000000000,-106.38,-12.845,-11.215,-15347.,-17935.
18.00000000000,-106.35,-12.846,-11.215,-15348.,-17937.
19.00000000000,-106.33,-12.848,-11.215,-15349.,-17940.
20.00000000000,-106.31,-12.849,-11.215,-15350.,-17942.
21.00000000000,-106.29,-12.851,-11.216,-15351.,-17944.
22.00000000000,-106.27,-12.853,-11.216,-15352.,-17946.
23.00000000000,-106.26,-12.855,-11.217,-15353.,-17947.
24.00000000000,-106.24,-12.856,-11.217,-15354.,-17949.
25.00000000000,-106.23,-12.858,-11.218,-15355.,-17950.
26.00000000000,-106.22,-12.860,-11.219,-15355.,-17952.
27.00000000000,-106.21,-12.862,-11.219,-15356.,-17953.
28.00000000000,-106.20,-12.863,-11.220,-15357.,-17954.
29.00000000000,-106.19,-12.865,-11.220,-15357.,-17955.
30.00000000000,-106.18,-12.866,-11.221,-15358.,-17957.
31.00000000000,-106.17,-12.868,-11.221,-15359.,-17958.
32.00000000000,-106.16,-12.870,-11.221,-15359.,-17959.
33.00000000000,-106.15,-12.871,-11.222,-15360.,-17960.
34.00000000000,-106.14,-12.873,-11.222,-15360.,-17961.
35.00000000000,-106.13,-12.874,-11.223,-15360.,-17962.
36.00000000000,-106.12,-12.875,-11.223,-15361.,-17963.
37.00000000000,-106.11,-12.877,-11.223,-15361.,-17964.
38.00000000000,-106.11,-12.878,-11.223,-15362.,-17964.
39.00000000000,-106.10,-12.879,-11.224,-15362.,-17965.
40.00000000000,-106.09,-12.881,-11.224,-15362.,-17966.
41.00000000000,-106.08,-12.882,-11.225,-15363.,-17966.
42.00000000000,-106.07,-12.883,-11.225,-15363.,-17967.
43.00000000000,-106.06,-12.884,-11.225,-15363.,-17967.
44.00000000000,-106.06,-12.885,-11.225,-15364.,-17968.
45.00000000000,-106.05,-12.886,-11.225,-15364.,-17968.
46.00000000000,-106.04,-12.887,-11.225,-15364.,-17969.
47.00000000000,-106.03,-12.888,-11.225,-15364.,-17969.
48.00000000000,-106.02,-12.889,-11.225,-15365.,-17970.
49.00000000000,-106.01,-12.889,-11.225,-15365.,-17970.
50.00000000000,-106.00,-12.890,-11.225,-15365.,-17971.
51.00000000000,-106.00,-12.891,-11.226,-15365.,-17971.
52.00000000000,-106.02,-12.897,-11.230,-15366.,-17971.
53.00000000000,-106.00,-12.896,-11.229,-15366.,-17972.
54.00000000000,-105.99,-12.896,-11.228,-15366.,-17972.
55.00000000000,-105.98,-12.896,-11.227,-15366.,-17972.
56.00000000000,-106.00,-12.901,-11.231,-15366.,-17973.
57.00000000000,-105.98,-12.900,-11.230,-15367.,-17973.
58.00000000000,-105.96,-12.900,-11.229,-15367.,-17973.
59.00000000000,-105.95,-12.900,-11.228,-15367.,-17973.
60.00000000000,-105.94,-12.900,-11.228,-15367.,-17974.
61.00000000000,-105.93,-12.901,-11.228,-15367.,-17974.
62.00000000000,-105.92,-12.901,-11.228,-15367.,-17974.
63.00000000000,-105.91,-12.902,-11.227,-15367.,-17975.
64.00000000000,-105.90,-12.903,-11.227,-15368.,-17975.
65.00000000000,-105.90,-12.903,-11.227,-15368.,-17975.
66.00000000000,-105.89,-12.904,-11.227,-15368.,-17975.
67.00000000000,-105.88,-12.905,-11.228,-15368.,-17976.
68.00000000000,-105.87,-12.906,-11.228,-15368.,-17976.
69.00000000000,-105.97,-12.919,-11.240,-15368.,-17976.
70.00000000000,-105.92,-12.916,-11.236,-15368.,-17976.
71.00000000000,-105.89,-12.914,-11.233,-15369.,-17977.
72.00000000000,-105.88,-12.913,-11.232,-15369.,-17977.
73.00000000000,-105.86,-12.912,-11.231,-15369.,-17977.
74.00000000000,-105.85,-12.912,-11.230,-15369.,-17977.
75.00000000000,-105.84,-12.913,-11.230,-15369.,-17977.
76.00000000000,-105.83,-12.913,-11.230,-15369.,-17978.
77.00000000000,-105.82,-12.914,-11.230,-15369.,-17978.
78.00000000000,-105.81,-12.914,-11.230,-15369.,-17978.
79.00000000000,-105.80,-12.915,-11.230,-15369.,-17978.
80.00000000000,-105.80,-12.916,-11.230,-15369.,-17978.
81.00000000000,-105.79,-12.916,-11.230,-15370.,-17979.
82.00000000000,-105.84,-12.925,-11.237,-15370.,-17979.
83.00000000000,-105.81,-12.923,-11.235,-15370.,-17979.
84.00000000000,-105.79,-12.922,-11.233,-15370.,-17979.
85.00000000000,-105.78,-12.922,-11.232,-15370.,-17979.
86.00000000000,-105.77,-12.922,-11.232,-15370.,-17979.
87.00000000000,-105.76,-12.922,-11.231,-15370.,-17980.
88.00000000000,-105.75,-12.922,-11.231,-15370.,-17980.
89.00000000000,-105.74,-12.923,-11.231,-15370.,-17980.
90.00000000000,-105.73,-12.923,-11.231,-15370.,-17980.
91.00000000000,-105.72,-12.924,-11.231,-15370.,-17980.
92.00000000000,-105.71,-12.925,-11.231,-15370.,-17980.
93.00000000000,-105.97,-12.957,-11.262,-15370.,-17981.
94.00000000000,-105.85,-12.947,-11.252,-15371.,-17981.
95.00000000000,-105.81,-12.940,-11.244,-15371.,-17981.
96.00000000000,-105.78,-12.937,-11.240,-15371.,-17981.
97.00000000000,-105.76,-12.935,-11.238,-15371.,-17981.
98.00000000000,-105.74,-12.934,-11.237,-15371.,-17981.
99.00000000000,-105.73,-12.933,-11.236,-15371.,-17981.
100.0000000000,-105.71,-12.933,-11.235,-15371.,-17981.
101.0000000000,-105.70,-12.933,-11.235,-15371.,-17982.
102.0000000000,-105.69,-12.934,-11.235,-15371.,-17982.
103.0000000000,-105.68,-12.934,-11.235,-15371.,-17982.
104.0000000000,-105.67,-12.935,-11.234,-15371.,-17982.
105.0000000000,-105.66,-12.935,-11.234,-15371.,-17982.
106.0000000000,-105.65,-12.936,-11.234,-15371.,-17982.
107.0000000000,-105.64,-12.936,-11.234,-15371.,-17982.
108.0000000000,-105.79,-12.955,-11.252,-15371.,-17982.
109.0000000000,-105.71,-12.949,-11.246,-15371.,-17982.
110.0000000000,-105.69,-12.946,-11.242,-15371.,-17983.
111.0000000000,-105.67,-12.944,-11.239,-15371.,-17983.
112.0000000000,-105.65,-12.943,-11.238,-15371.,-17983.
113.0000000000,-105.64,-12.942,-11.237,-15371.,-17983.
114.0000000000,-105.63,-12.942,-11.237,-15371.,-17983.
115.0000000000,-105.62,-12.942,-11.236,-15371.,-17983.
116.0000000000,-105.61,-12.942,-11.236,-15372.,-17983.
117.0000000000,-105.60,-12.943,-11.236,-15372.,-17983.
118.0000000000,-106.09,-13.001,-11.294,-15372.,-17983.
119.0000000000,-106.72,-13.079,-11.372,-15372.,-17983.
120.0000000000,-106.27,-13.033,-11.325,-15372.,-17984.
121.0000000000,-106.11,-13.005,-11.295,-15372.,-17984.
122.0000000000,-106.34,-13.025,-11.316,-15372.,-17984.
123.0000000000,-106.13,-13.001,-11.294,-15373.,-17984.
124.0000000000,-106.03,-12.986,-11.279,-15373.,-17984.
125.0000000000,-105.97,-12.977,-11.271,-15373.,-17984.
126.0000000000,-105.92,-12.971,-11.266,-15373.,-17984.
127.0000000000,-105.88,-12.968,-11.263,-15373.,-17984.
128.0000000000,-105.85,-12.966,-11.261,-15373.,-17984.
129.0000000000,-105.82,-12.964,-11.259,-15373.,-17984.
130.0000000000,-105.96,-12.983,-11.277,-15373.,-17984.
131.0000000000,-106.07,-12.999,-11.293,-15373.,-17984.
132.0000000000,-105.94,-12.987,-11.281,-15373.,-17984.
133.0000000000,-105.89,-12.979,-11.272,-15373.,-17984.
134.0000000000,-105.85,-12.974,-11.268,-15373.,-17984.
135.0000000000,-106.09,-13.003,-11.296,-15373.,-17984.
136.0000000000,-105.95,-12.990,-11.284,-15373.,-17984.
137.0000000000,-105.90,-12.982,-11.275,-15373.,-17984.
138.0000000000,-105.86,-12.977,-11.271,-15373.,-17984.
139.0000000000,-105.83,-12.975,-11.268,-15373.,-17984.
140.0000000000,-105.81,-12.973,-11.266,-15374.,-17984.
141.0000000000,-105.79,-12.972,-11.265,-15374.,-17984.
142.0000000000,-105.77,-12.971,-11.264,-15374.,-17984.
143.0000000000,-105.76,-12.971,-11.264,-15374.,-17984.
144.0000000000,-106.35,-13.040,-11.332,-15374.,-17984.
145.0000000000,-106.12,-13.022,-11.314,-15374.,-17984.
146.0000000000,-106.94,-13.113,-11.403,-15374.,-17985.
147.0000000000,-106.47,-13.064,-11.356,-15375.,-17985.
148.0000000000,-106.30,-13.035,-11.326,-15375.,-17985.
149.0000000000,-106.33,-13.033,-11.324,-15375.,-17985.
150.0000000000,-106.20,-13.016,-11.309,-15375.,-17985.
151.0000000000,-106.12,-13.006,-11.299,-15375.,-17985.
152.0000000000,-106.07,-12.999,-11.294,-15375.,-17985.
153.0000000000,-106.03,-12.995,-11.290,-15375.,-17985.
154.0000000000,-106.01,-12.995,-11.290,-15375.,-17985.
155.0000000000,-105.97,-12.992,-11.288,-15375.,-17985.
156.0000000000,-105.94,-12.991,-11.286,-15375.,-17985.
157.0000000000,-105.92,-12.990,-11.285,-15375.,-17985.
158.0000000000,-105.91,-12.989,-11.284,-15375.,-17985.
159.0000000000,-106.10,-13.014,-11.308,-15375.,-17985.
160.0000000000,-105.99,-13.005,-11.299,-15375.,-17985.
161.0000000000,-105.95,-12.999,-11.293,-15375.,-17985.
162.0000000000,-105.92,-12.996,-11.290,-15376.,-17985.
163.0000000000,-105.90,-12.994,-11.287,-15376.,-17985.
164.0000000000,-105.88,-12.992,-11.286,-15376.,-17985.
165.0000000000,-106.00,-13.008,-11.301,-15376.,-17985.
166.0000000000,-107.13,-13.139,-11.433,-15376.,-17986.
167.0000000000,-106.65,-13.098,-11.392,-15376.,-17986.
168.0000000000,-106.43,-13.063,-11.354,-15376.,-17986.
169.0000000000,-106.40,-13.052,-11.344,-15377.,-17986.
170.0000000000,-106.31,-13.038,-11.331,-15377.,-17986.
171.0000000000,-106.23,-13.026,-11.321,-15377.,-17986.
172.0000000000,-106.17,-13.018,-11.314,-15377.,-17986.
173.0000000000,-106.12,-13.013,-11.310,-15377.,-17986.
174.0000000000,-106.08,-13.010,-11.307,-15377.,-17986.
175.0000000000,-106.05,-13.008,-11.305,-15377.,-17986.
176.0000000000,-106.03,-13.007,-11.304,-15377.,-17986.
177.0000000000,-106.00,-13.006,-11.303,-15377.,-17986.
178.0000000000,-105.98,-13.005,-11.302,-15377.,-17986.
179.0000000000,-105.97,-13.005,-11.301,-15377.,-17986.
180.0000000000,-105.95,-13.004,-11.301,-15377.,-17986.
181.0000000000,-106.24,-13.039,-11.335,-15377.,-17986.
182.0000000000,-106.10,-13.027,-11.323,-15377.,-17986.
183.0000000000,-106.11,-13.028,-11.322,-15377.,-17986.
184.0000000000,-106.05,-13.020,-11.315,-15378.,-17986.
185.0000000000,-106.01,-13.015,-11.311,-15378.,-17987.
186.0000000000,-105.99,-13.012,-11.308,-15378.,-17987.
187.0000000000,-105.96,-13.011,-11.306,-15378.,-17987.
188.0000000000,-105.94,-13.009,-11.305,-15378.,-17987.
189.0000000000,-105.93,-13.009,-11.304,-15378.,-17987.
190.0000000000,-105.91,-13.008,-11.303,-15378.,-17987.
191.0000000000,-105.90,-13.008,-11.303,-15378.,-17987.
192.0000000000,-105.89,-13.007,-11.302,-15378.,-17987.
193.0000000000,-105.88,-13.007,-11.302,-15378.,-17987.
194.0000000000,-105.86,-13.007,-11.301,-15378.,-17987.
195.0000000000,-105.85,-13.007,-11.301,-15378.,-17987.
196.0000000000,-105.92,-13.017,-11.310,-15378.,-17987.
197.0000000000,-106.66,-13.103,-11.396,-15379.,-17987.
198.0000000000,-106.71,-13.117,-11.411,-15379.,-17987.
199.0000000000,-106.49,-13.090,-11.382,-15379.,-17988.
200.0000000000,-106.45,-13.079,-11.370,-15379.,-17988.
201.0000000000,-106.31,-13.057,-11.350,-15379.,-17988.
202.0000000000,-106.25,-13.047,-11.340,-15379.,-17988.
203.0000000000,-106.21,-13.042,-11.336,-15380.,-17988.
204.0000000000,-106.15,-13.034,-11.330,-15380.,-17988.
205.0000000000,-106.11,-13.029,-11.326,-15380.,-17988.
206.0000000000,-106.07,-13.026,-11.323,-15380.,-17988.
207.0000000000,-106.04,-13.023,-11.321,-15380.,-17988.
208.0000000000,-106.05,-13.027,-11.324,-15380.,-17988.
209.0000000000,-106.02,-13.024,-11.321,-15380.,-17988.
210.0000000000,-106.11,-13.036,-11.333,-15380.,-17988.
211.0000000000,-106.04,-13.030,-11.327,-15380.,-17988.
212.0000000000,-106.01,-13.026,-11.323,-15380.,-17988.
213.0000000000,-105.98,-13.024,-11.321,-15380.,-17988.
214.0000000000,-105.97,-13.022,-11.320,-15380.,-17988.
215.0000000000,-105.95,-13.021,-11.318,-15380.,-17988.
216.0000000000,-105.93,-13.020,-11.318,-15380.,-17988.
217.0000000000,-105.92,-13.020,-11.317,-15380.,-17988.
218.0000000000,-105.91,-13.020,-11.316,-15380.,-17988.
219.0000000000,-105.90,-13.019,-11.316,-15380.,-17988.
220.0000000000,-105.88,-13.019,-11.315,-15380.,-17988.
221.0000000000,-105.87,-13.019,-11.315,-15381.,-17988.
222.0000000000,-105.86,-13.019,-11.315,-15381.,-17988.
223.0000000000,-105.86,-13.019,-11.315,-15381.,-17988.
224.0000000000,-105.89,-13.024,-11.319,-15381.,-17988.
225.0000000000,-105.86,-13.022,-11.317,-15381.,-17988.
226.0000000000,-105.84,-13.020,-11.316,-15381.,-17988.
227.0000000000,-105.83,-13.019,-11.315,-15381.,-17988.
228.0000000000,-105.82,-13.019,-11.314,-15381.,-17988.
229.0000000000,-105.81,-13.018,-11.314,-15381.,-17988.
230.0000000000,-105.80,-13.018,-11.313,-15381.,-17988.
231.0000000000,-105.79,-13.018,-11.313,-15381.,-17988.
232.0000000000,-105.78,-13.018,-11.312,-15381.,-17988.
233.0000000000,-105.77,-13.017,-11.312,-15381.,-17988.
234.0000000000,-105.79,-13.021,-11.315,-15381.,-17988.
235.0000000000,-105.77,-13.019,-11.313,-15381.,-17988.
236.0000000000,-106.39,-13.091,-11.384,-15382.,-17989.
237.0000000000,-106.11,-13.067,-11.361,-15382.,-17989.
238.0000000000,-106.10,-13.061,-11.354,-15382.,-17989.
239.0000000000,-106.82,-13.140,-11.433,-15382.,-17989.
240.0000000000,-107.07,-13.174,-11.469,-15382.,-17990.
241.0000000000,-106.63,-13.122,-11.417,-15383.,-17990.
242.0000000000,-106.45,-13.090,-11.384,-15383.,-17990.
243.0000000000,-106.34,-13.069,-11.366,-15383.,-17990.
244.0000000000,-106.26,-13.057,-11.356,-15383.,-17990.
245.0000000000,-106.19,-13.049,-11.349,-15383.,-17990.
246.0000000000,-106.43,-13.077,-11.377,-15383.,-17990.
247.0000000000,-106.26,-13.061,-11.363,-15383.,-17989.
248.0000000000,-106.41,-13.078,-11.379,-15383.,-17989.
249.0000000000,-106.40,-13.079,-11.381,-15383.,-17990.
250.0000000000,-106.27,-13.063,-11.366,-15383.,-17990.
251.0000000000,-106.21,-13.054,-11.357,-15383.,-17990.
252.0000000000,-106.34,-13.069,-11.372,-15383.,-17990.
253.0000000000,-106.26,-13.062,-11.365,-15383.,-17990.
254.0000000000,-106.28,-13.064,-11.367,-15383.,-17990.
255.0000000000,-106.20,-13.054,-11.359,-15383.,-17990.
256.0000000000,-106.15,-13.048,-11.353,-15383.,-17990.
257.0000000000,-106.12,-13.045,-11.350,-15383.,-17990.
258.0000000000,-106.09,-13.042,-11.347,-15383.,-17989.
259.0000000000,-106.07,-13.040,-11.346,-15383.,-17989.
260.0000000000,-106.20,-13.057,-11.362,-15383.,-17989.
261.0000000000,-106.42,-13.085,-11.390,-15383.,-17989.
262.0000000000,-106.32,-13.076,-11.382,-15383.,-17990.
263.0000000000,-108.01,-13.267,-11.573,-15384.,-17990.
264.0000000000,-108.62,-13.352,-11.661,-15384.,-17991.
265.0000000000,-107.69,-13.245,-11.552,-15385.,-17992.
266.0000000000,-107.34,-13.180,-11.485,-15385.,-17992.
267.0000000000,-107.13,-13.138,-11.447,-15385.,-17992.
268.0000000000,-106.97,-13.112,-11.426,-15385.,-17992.
269.0000000000,-106.85,-13.096,-11.412,-15385.,-17992.
270.0000000000,-106.76,-13.085,-11.404,-15385.,-17992.
271.0000000000,-106.69,-13.078,-11.398,-15385.,-17991.
272.0000000000,-106.87,-13.102,-11.422,-15385.,-17991.
273.0000000000,-106.71,-13.088,-11.410,-15385.,-17991.
274.0000000000,-106.64,-13.080,-11.401,-15385.,-17991.
275.0000000000,-106.59,-13.074,-11.396,-15384.,-17990.
276.0000000000,-106.55,-13.071,-11.393,-15384.,-17990.
277.0000000000,-106.51,-13.068,-11.390,-15384.,-17990.
278.0000000000,-106.48,-13.066,-11.389,-15384.,-17990.
279.0000000000,-106.46,-13.065,-11.388,-15384.,-17990.
280.0000000000,-106.44,-13.064,-11.386,-15384.,-17990.
281.0000000000,-106.42,-13.063,-11.385,-15384.,-17990.
282.0000000000,-106.40,-13.062,-11.384,-15384.,-17990.
283.0000000000,-106.38,-13.062,-11.384,-15385.,-17990.
284.0000000000,-106.37,-13.061,-11.383,-15385.,-17990.
285.0000000000,-106.36,-13.061,-11.382,-15385.,-17990.
286.0000000000,-106.35,-13.061,-11.382,-15385.,-17990.
287.0000000000,-106.55,-13.086,-11.407,-15385.,-17990.
288.0000000000,-106.84,-13.122,-11.443,-15385.,-17990.
289.0000000000,-107.83,-13.238,-11.559,-15385.,-17990.
290.0000000000,-107.25,-13.180,-11.501,-15385.,-17991.
291.0000000000,-107.02,-13.141,-11.460,-15385.,-17991.
292.0000000000,-106.90,-13.117,-11.438,-15386.,-17991.
293.0000000000,-106.81,-13.101,-11.424,-15385.,-17991.
294.0000000000,-106.73,-13.091,-11.416,-15385.,-17991.
295.0000000000,-106.68,-13.084,-11.410,-15385.,-17990.
296.0000000000,-106.63,-13.080,-11.407,-15385.,-17990.
297.0000000000,-106.59,-13.077,-11.404,-15385.,-17990.
298.0000000000,-106.56,-13.075,-11.402,-15385.,-17990.
299.0000000000,-106.53,-13.073,-11.401,-15385.,-17990.
300.0000000000,-106.51,-13.072,-11.399,-15385.,-17990.
301.0000000000,-106.49,-13.071,-11.398,-15385.,-17990.
302.0000000000,-106.47,-13.070,-11.397,-15385.,-17990.
303.0000000000,-106.45,-13.069,-11.397,-15385.,-17990.
304.0000000000,-106.45,-13.070,-11.397,-15385.,-17990.
305.0000000000,-106.43,-13.069,-11.396,-15385.,-17990.
306.0000000000,-106.41,-13.068,-11.395,-15386.,-17990.
307.0000000000,-106.40,-13.067,-11.394,-15386.,-17990.
308.0000000000,-106.55,-13.085,-11.411,-15386.,-17990.
309.0000000000,-106.51,-13.084,-11.410,-15386.,-17990.
310.0000000000,-106.59,-13.093,-11.419,-15386.,-17990.
311.0000000000,-106.61,-13.097,-11.422,-15386.,-17990.
312.0000000000,-106.52,-13.086,-11.412,-15386.,-17990.
313.0000000000,-106.61,-13.094,-11.420,-15386.,-17990.
314.0000000000,-106.52,-13.084,-11.411,-15386.,-17990.
315.0000000000,-106.48,-13.078,-11.405,-15386.,-17990.
316.0000000000,-106.48,-13.078,-11.404,-15386.,-17990.
317.0000000000,-106.45,-13.075,-11.402,-15386.,-17990.
318.0000000000,-106.42,-13.072,-11.399,-15386.,-17990.
319.0000000000,-106.40,-13.070,-11.397,-15386.,-17990.
320.0000000000,-106.38,-13.068,-11.395,-15386.,-17990.
321.0000000000,-106.36,-13.067,-11.394,-15386.,-17990.
322.0000000000,-106.35,-13.066,-11.393,-15386.,-17990.
323.0000000000,-106.33,-13.065,-11.392,-15386.,-17990.
324.0000000000,-106.32,-13.064,-11.392,-15386.,-17989.
325.0000000000,-106.31,-13.064,-11.391,-15386.,-17989.
326.0000000000,-106.35,-13.069,-11.396,-15386.,-17989.
327.0000000000,-106.36,-13.073,-11.399,-15386.,-17989.
328.0000000000,-106.65,-13.106,-11.432,-15386.,-17990.
329.0000000000,-106.75,-13.121,-11.447,-15386.,-17990.
330.0000000000,-106.58,-13.101,-11.427,-15386.,-17990.
331.0000000000,-106.50,-13.088,-11.414,-15386.,-17990.
332.0000000000,-106.45,-13.080,-11.407,-15386.,-17990.
333.0000000000,-106.42,-13.074,-11.402,-15387.,-17990.
334.0000000000,-106.39,-13.071,-11.399,-15387.,-17990.
335.0000000000,-106.36,-13.068,-11.397,-15386.,-17989.
336.0000000000,-106.34,-13.066,-11.395,-15386.,-17989.
337.0000000000,-106.32,-13.065,-11.394,-15386.,-17989.
338.0000000000,-106.31,-13.064,-11.393,-15386.,-17989.
339.0000000000,-106.29,-13.063,-11.392,-15387.,-17989.
340.0000000000,-106.34,-13.070,-11.398,-15387.,-17989.
341.0000000000,-106.30,-13.067,-11.395,-15387.,-17989.
342.0000000000,-106.28,-13.064,-11.393,-15387.,-17989.
343.0000000000,-106.26,-13.063,-11.391,-15387.,-17989.
344.0000000000,-106.25,-13.061,-11.390,-15387.,-17989.
345.0000000000,-106.24,-13.060,-11.389,-15387.,-17989.
346.0000000000,-106.22,-13.060,-11.388,-15387.,-17989.
347.0000000000,-106.21,-13.059,-11.387,-15387.,-17989.
348.0000000000,-106.20,-13.058,-11.387,-15387.,-17989.
349.0000000000,-106.19,-13.058,-11.386,-15387.,-17989.
350.0000000000,-106.18,-13.057,-11.385,-15387.,-17989.
351.0000000000,-106.17,-13.056,-11.385,-15387.,-17989.
352.0000000000,-106.16,-13.056,-11.384,-15387.,-17989.
353.0000000000,-106.15,-13.055,-11.383,-15387.,-17989.
354.0000000000,-106.14,-13.055,-11.383,-15387.,-17989.
355.0000000000,-106.37,-13.082,-11.410,-15387.,-17989.
356.0000000000,-106.35,-13.083,-11.410,-15387.,-17989.
357.0000000000,-106.27,-13.073,-11.400,-15387.,-17989.
358.0000000000,-106.23,-13.066,-11.393,-15387.,-17989.
359.0000000000,-106.20,-13.062,-11.390,-15387.,-17989.
360.0000000000,-106.26,-13.069,-11.396,-15387.,-17989.
361.0000000000,-106.37,-13.082,-11.410,-15387.,-17989.
362.0000000000,-106.41,-13.088,-11.416,-15387.,-17989.
363.0000000000,-106.31,-13.076,-11.404,-15387.,-17989.
364.0000000000,-106.26,-13.068,-11.397,-15387.,-17989.
365.0000000000,-106.23,-13.063,-11.392,-15387.,-17989.
366.0000000000,-106.20,-13.060,-11.389,-15387.,-17989.
367.0000000000,-106.18,-13.058,-11.387,-15387.,-17989.
368.0000000000,-106.16,-13.056,-11.386,-15387.,-17989.
369.0000000000,-106.14,-13.054,-11.384,-15387.,-17988.
370.0000000000,-106.13,-13.053,-11.383,-15387.,-17988.
371.0000000000,-106.11,-13.052,-11.383,-15387.,-17988.
372.0000000000,-106.10,-13.052,-11.382,-15387.,-17988.
373.0000000000,-106.09,-13.051,-11.381,-15387.,-17988.
374.0000000000,-106.08,-13.050,-11.380,-15387.,-17988.
375.0000000000,-106.07,-13.050,-11.380,-15387.,-17988.
376.0000000000,-106.06,-13.049,-11.379,-15387.,-17988.
377.0000000000,-106.05,-13.048,-11.378,-15387.,-17988.
378.0000000000,-106.04,-13.048,-11.378,-15387.,-17988.
379.0000000000,-106.03,-13.047,-11.377,-15387.,-17988.
380.0000000000,-106.02,-13.047,-11.376,-15387.,-17988.
381.0000000000,-106.01,-13.046,-11.376,-15387.,-17988.
382.0000000000,-106.00,-13.046,-11.375,-15388.,-17988.
383.0000000000,-105.99,-13.045,-11.375,-15388.,-17988.
384.0000000000,-105.99,-13.044,-11.374,-15388.,-17988.
385.0000000000,-105.98,-13.044,-11.374,-15388.,-17988.
386.0000000000,-105.97,-13.043,-11.373,-15388.,-17988.
387.0000000000,-105.96,-13.043,-11.372,-15388.,-17988.
388.0000000000,-105.95,-13.042,-11.372,-15388.,-17988.
389.0000000000,-105.96,-13.045,-11.374,-15388.,-17988.
390.0000000000,-105.95,-13.043,-11.372,-15388.,-17988.
391.0000000000,-105.94,-13.042,-11.371,-15388.,-17988.
392.0000000000,-105.93,-13.041,-11.370,-15388.,-17988.
393.0000000000,-105.92,-13.040,-11.370,-15388.,-17987.
394.0000000000,-105.91,-13.040,-11.369,-15388.,-17987.
395.0000000000,-105.90,-13.039,-11.368,-15388.,-17987.
396.0000000000,-105.89,-13.038,-11.368,-15388.,-17987.
397.0000000000,-105.88,-13.038,-11.367,-15388.,-17987.
398.0000000000,-105.87,-13.037,-11.366,-15388.,-17987.
399.0000000000,-105.87,-13.037,-11.366,-15388.,-17987.
400.0000000000,-105.86,-13.036,-11.365,-15388.,-17987.
401.0000000000,-105.85,-13.036,-11.365,-15388.,-17987.
402.0000000000,-105.84,-13.035,-11.364,-15388.,-17987.
403.0000000000,-105.83,-13.035,-11.364,-15388.,-17987.
404.0000000000,-105.82,-13.034,-11.363,-15388.,-17987.
405.0000000000,-105.82,-13.033,-11.362,-15388.,-17987.
406.0000000000,-105.81,-13.033,-11.362,-15388.,-17987.
407.0000000000,-105.80,-13.032,-11.361,-15388.,-17987.
408.0000000000,-105.79,-13.032,-11.361,-15388.,-17987.
409.0000000000,-105.78,-13.031,-11.360,-15388.,-17987.
410.0000000000,-105.78,-13.031,-11.360,-15388.,-17987.
411.0000000000,-105.77,-13.030,-11.359,-15388.,-17987.
412.0000000000,-105.76,-13.030,-11.359,-15388.,-17987.
413.0000000000,-105.75,-13.029,-11.358,-15388.,-17987.
414.0000000000,-105.75,-13.029,-11.358,-15388.,-17987.
415.0000000000,-105.74,-13.028,-11.357,-15388.,-17987.
416.0000000000,-105.73,-13.028,-11.356,-15388.,-17987.
417.0000000000,-105.72,-13.027,-11.356,-15388.,-17987.
418.0000000000,-105.71,-13.027,-11.355,-15388.,-17986.
419.0000000000,-105.71,-13.026,-11.355,-15388.,-17986.
420.0000000000,-105.70,-13.026,-11.354,-15388.,-17986.
421.0000000000,-105.71,-13.027,-11.356,-15388.,-17986.
422.0000000000,-105.90,-13.051,-11.378,-15388.,-17986.
423.0000000000,-105.86,-13.049,-11.377,-15388.,-17986.
424.0000000000,-105.80,-13.040,-11.368,-15388.,-17987.
425.0000000000,-105.77,-13.035,-11.363,-15388.,-17986.
426.0000000000,-105.75,-13.032,-11.360,-15388.,-17986.
427.0000000000,-105.73,-13.029,-11.358,-15388.,-17986.
428.0000000000,-105.71,-13.027,-11.356,-15388.,-17986.
429.0000000000,-105.70,-13.025,-11.355,-15388.,-17986.
430.0000000000,-105.69,-13.024,-11.354,-15388.,-17986.
431.0000000000,-105.68,-13.023,-11.353,-15388.,-17986.
432.0000000000,-105.66,-13.022,-11.352,-15388.,-17986.
433.0000000000,-105.65,-13.022,-11.351,-15388.,-17986.
434.0000000000,-105.65,-13.023,-11.352,-15388.,-17986.
435.0000000000,-105.64,-13.022,-11.351,-15388.,-17986.
436.0000000000,-105.63,-13.021,-11.350,-15388.,-17986.
437.0000000000,-105.62,-13.020,-11.350,-15388.,-17986.
438.0000000000,-105.61,-13.019,-11.349,-15388.,-17986.
439.0000000000,-105.61,-13.019,-11.348,-15388.,-17986.
440.0000000000,-105.60,-13.018,-11.348,-15388.,-17986.
441.0000000000,-105.59,-13.017,-11.347,-15388.,-17986.
442.0000000000,-105.58,-13.017,-11.347,-15388.,-17986.
443.0000000000,-105.57,-13.016,-11.346,-15388.,-17986.
444.0000000000,-105.57,-13.016,-11.345,-15388.,-17986.
445.0000000000,-105.56,-13.015,-11.345,-15388.,-17986.
446.0000000000,-105.55,-13.015,-11.344,-15388.,-17986.
447.0000000000,-105.54,-13.014,-11.344,-15388.,-17986.
448.0000000000,-105.58,-13.020,-11.349,-15388.,-17986.
449.0000000000,-105.55,-13.017,-11.347,-15388.,-17986.
450.0000000000,-105.54,-13.016,-11.345,-15388.,-17986.
451.0000000000,-105.54,-13.016,-11.345,-15388.,-17986.
452.0000000000,-105.52,-13.014,-11.343,-15388.,-17985.
453.0000000000,-105.51,-13.013,-11.342,-15388.,-17985.
454.0000000000,-105.51,-13.012,-11.342,-15388.,-17985.
455.0000000000,-105.50,-13.011,-11.341,-15388.,-17985.
456.0000000000,-105.49,-13.011,-11.340,-15388.,-17985.
457.0000000000,-105.48,-13.010,-11.340,-15388.,-17985.
458.0000000000,-105.47,-13.010,-11.339,-15388.,-17985.
459.0000000000,-105.64,-13.030,-11.359,-15388.,-17985.
460.0000000000,-105.56,-13.022,-11.351,-15388.,-17985.
461.0000000000,-105.53,-13.019,-11.347,-15388.,-17985.
462.0000000000,-105.51,-13.015,-11.344,-15388.,-17985.
463.0000000000,-105.51,-13.015,-11.344,-15388.,-17985.
464.0000000000,-105.49,-13.013,-11.342,-15388.,-17985.
465.0000000000,-105.47,-13.011,-11.340,-15388.,-17985.
466.0000000000,-105.46,-13.009,-11.339,-15388.,-17985.
467.0000000000,-105.45,-13.008,-11.338,-15388.,-17985.
468.0000000000,-105.44,-13.007,-11.337,-15388.,-17985.
469.0000000000,-105.43,-13.007,-11.337,-15388.,-17985.
470.0000000000,-105.42,-13.006,-11.336,-15388.,-17985.
471.0000000000,-105.41,-13.005,-11.335,-15388.,-17985.
472.0000000000,-105.40,-13.004,-11.335,-15388.,-17985.
473.0000000000,-105.40,-13.004,-11.334,-15388.,-17985.
474.0000000000,-105.39,-13.003,-11.333,-15388.,-17985.
475.0000000000,-105.40,-13.006,-11.336,-15388.,-17985.
476.0000000000,-105.39,-13.005,-11.334,-15388.,-17985.
477.0000000000,-105.38,-13.003,-11.333,-15388.,-17984.
478.0000000000,-105.37,-13.002,-11.332,-15388.,-17984.
479.0000000000,-105.36,-13.002,-11.331,-15388.,-17984.
480.0000000000,-105.35,-13.001,-11.331,-15388.,-17984.
481.0000000000,-105.34,-13.000,-11.330,-15388.,-17984.
482.0000000000,-105.33,-13.000,-11.330,-15388.,-17984.
483.0000000000,-105.33,-12.999,-11.329,-15388.,-17984.
484.0000000000,-105.32,-12.999,-11.329,-15388.,-17984.
485.0000000000,-105.31,-12.998,-11.328,-15388.,-17984.
486.0000000000,-105.30,-12.998,-11.328,-15388.,-17984.
487.0000000000,-105.30,-12.997,-11.327,-15388.,-17984.
488.0000000000,-105.29,-12.997,-11.327,-15388.,-17984.
489.0000000000,-105.28,-12.996,-11.326,-15388.,-17984.
490.0000000000,-105.28,-12.996,-11.325,-15388.,-17984.
491.0000000000,-105.27,-12.995,-11.325,-15388.,-17984.
492.0000000000,-105.40,-13.011,-11.340,-15388.,-17984.
493.0000000000,-105.33,-13.005,-11.334,-15388.,-17984.
494.0000000000,-105.37,-13.008,-11.337,-15388.,-17984.
495.0000000000,-105.44,-13.017,-11.346,-15388.,-17984.
496.0000000000,-105.37,-13.009,-11.338,-15388.,-17984.
497.0000000000,-105.34,-13.004,-11.334,-15388.,-17984.
498.0000000000,-105.45,-13.016,-11.345,-15388.,-17984.
499.0000000000,-105.40,-13.012,-11.342,-15388.,-17984.
500.0000000000,-105.35,-13.006,-11.335,-15388.,-17984.
501.0000000000,-105.33,-13.002,-11.332,-15388.,-17984.
502.0000000000,-105.31,-12.999,-11.329,-15388.,-17984.
503.0000000000,-105.29,-12.997,-11.327,-15388.,-17983.
504.0000000000,-105.28,-12.995,-11.326,-15388.,-17983.
505.0000000000,-105.26,-12.994,-11.325,-15388.,-17983.
506.0000000000,-105.25,-12.993,-11.324,-15388.,-17983.
507.0000000000,-105.24,-12.992,-11.324,-15388.,-17983.
508.0000000000,-105.28,-12.998,-11.329,-15388.,-17983.
509.0000000000,-105.25,-12.995,-11.327,-15388.,-17983.
510.0000000000,-105.36,-13.009,-11.339,-15388.,-17983.
511.0000000000,-106.14,-13.098,-11.429,-15388.,-17983.
512.0000000000,-105.79,-13.067,-11.398,-15388.,-17983.
513.0000000000,-105.64,-13.041,-11.371,-15388.,-17984.
514.0000000000,-105.55,-13.025,-11.356,-15388.,-17983.
515.0000000000,-105.50,-13.014,-11.347,-15388.,-17983.
516.0000000000,-105.45,-13.008,-11.341,-15388.,-17983.
517.0000000000,-105.42,-13.003,-11.338,-15388.,-17983.
518.0000000000,-105.39,-13.000,-11.335,-15388.,-17983.
519.0000000000,-105.36,-12.998,-11.333,-15388.,-17983.
520.0000000000,-105.34,-12.997,-11.332,-15388.,-17983.
521.0000000000,-105.32,-12.995,-11.331,-15388.,-17983.
522.0000000000,-105.31,-12.994,-11.330,-15388.,-17982.
523.0000000000,-105.29,-12.993,-11.329,-15388.,-17982.
524.0000000000,-105.28,-12.992,-11.328,-15388.,-17982.
525.0000000000,-105.28,-12.994,-11.329,-15388.,-17982.
526.0000000000,-105.28,-12.994,-11.329,-15388.,-17982.
527.0000000000,-105.26,-12.993,-11.328,-15388.,-17982.
528.0000000000,-105.28,-12.995,-11.330,-15388.,-17982.
529.0000000000,-105.43,-13.013,-11.348,-15388.,-17982.
530.0000000000,-105.66,-13.042,-11.376,-15388.,-17982.
531.0000000000,-105.49,-13.023,-11.359,-15388.,-17982.
532.0000000000,-105.42,-13.012,-11.347,-15388.,-17982.
533.0000000000,-105.38,-13.004,-11.340,-15388.,-17982.
534.0000000000,-105.35,-12.999,-11.336,-15388.,-17982.
535.0000000000,-105.32,-12.996,-11.333,-15388.,-17982.
536.0000000000,-107.15,-13.204,-11.542,-15388.,-17982.
537.0000000000,-107.09,-13.217,-11.558,-15389.,-17983.
538.0000000000,-106.74,-13.171,-11.507,-15389.,-17983.
539.0000000000,-106.38,-13.112,-11.449,-15389.,-17983.
540.0000000000,-106.20,-13.078,-11.417,-15389.,-17983.
541.0000000000,-106.74,-13.131,-11.474,-15389.,-17983.
542.0000000000,-106.34,-13.089,-11.435,-15389.,-17983.
543.0000000000,-106.17,-13.063,-11.409,-15389.,-17983.
544.0000000000,-106.06,-13.047,-11.395,-15389.,-17983.
545.0000000000,-105.98,-13.036,-11.386,-15389.,-17983.
546.0000000000,-105.91,-13.028,-11.380,-15389.,-17982.
547.0000000000,-105.85,-13.023,-11.375,-15389.,-17982.
548.0000000000,-105.81,-13.020,-11.372,-15388.,-17982.
549.0000000000,-105.78,-13.017,-11.370,-15388.,-17981.
550.0000000000,-105.74,-13.015,-11.368,-15388.,-17981.
551.0000000000,-105.72,-13.013,-11.367,-15388.,-17981.
552.0000000000,-105.70,-13.012,-11.366,-15388.,-17981.
553.0000000000,-105.68,-13.011,-11.365,-15388.,-17981.
554.0000000000,-105.66,-13.010,-11.364,-15388.,-17981.
555.0000000000,-105.64,-13.009,-11.363,-15388.,-17980.
556.0000000000,-105.64,-13.010,-11.363,-15388.,-17980.
557.0000000000,-105.63,-13.011,-11.363,-15388.,-17980.
558.0000000000,-105.76,-13.026,-11.378,-15388.,-17980.
559.0000000000,-105.68,-13.019,-11.371,-15388.,-17980.
560.0000000000,-105.65,-13.014,-11.367,-15388.,-17980.
561.0000000000,-105.63,-13.011,-11.364,-15388.,-17980.
562.0000000000,-105.79,-13.031,-11.383,-15388.,-17980.
563.0000000000,-105.92,-13.047,-11.400,-15388.,-17980.
564.0000000000,-105.95,-13.052,-11.404,-15388.,-17980.
565.0000000000,-105.82,-13.035,-11.388,-15388.,-17980.
566.0000000000,-105.76,-13.025,-11.378,-15388.,-17980.
567.0000000000,-105.72,-13.019,-11.372,-15388.,-17980.
568.0000000000,-105.69,-13.014,-11.368,-15388.,-17979.
569.0000000000,-105.66,-13.011,-11.366,-15388.,-17979.
570.0000000000,-105.64,-13.009,-11.364,-15388.,-17979.
571.0000000000,-105.70,-13.017,-11.371,-15388.,-17979.
572.0000000000,-105.65,-13.013,-11.367,-15388.,-17979.
573.0000000000,-105.62,-13.010,-11.364,-15388.,-17979.
574.0000000000,-105.60,-13.007,-11.362,-15388.,-17979.
575.0000000000,-105.59,-13.006,-11.360,-15388.,-17979.
576.0000000000,-105.57,-13.004,-11.359,-15388.,-17979.
577.0000000000,-105.56,-13.003,-11.358,-15388.,-17979.
578.0000000000,-105.55,-13.003,-11.357,-15388.,-17978.
579.0000000000,-105.87,-13.040,-11.394,-15388.,-17978.
580.0000000000,-106.57,-13.124,-11.478,-15388.,-17979.
581.0000000000,-106.13,-13.080,-11.436,-15388.,-17979.
582.0000000000,-105.99,-13.054,-11.407,-15388.,-17979.
583.0000000000,-105.90,-13.037,-11.392,-15388.,-17979.
584.0000000000,-105.84,-13.027,-11.382,-15388.,-17979.
585.0000000000,-105.79,-13.020,-11.377,-15388.,-17979.
586.0000000000,-105.75,-13.015,-11.373,-15388.,-17978.
587.0000000000,-105.72,-13.012,-11.370,-15388.,-17978.
588.0000000000,-105.69,-13.010,-11.368,-15388.,-17978.
589.0000000000,-105.75,-13.019,-11.377,-15388.,-17978.
590.0000000000,-105.90,-13.038,-11.396,-15388.,-17978.
591.0000000000,-105.78,-13.026,-11.384,-15388.,-17978.
592.0000000000,-105.73,-13.018,-11.376,-15387.,-17978.
593.0000000000,-105.70,-13.013,-11.372,-15387.,-17978.
594.0000000000,-105.73,-13.016,-11.375,-15387.,-17977.
595.0000000000,-105.94,-13.042,-11.401,-15387.,-17978.
596.0000000000,-106.13,-13.066,-11.425,-15387.,-17978.
597.0000000000,-105.93,-13.044,-11.403,-15388.,-17978.
598.0000000000,-105.85,-13.030,-11.389,-15388.,-17978.
599.0000000000,-105.80,-13.021,-11.381,-15387.,-17977.
600.0000000000,-105.76,-13.016,-11.376,-15387.,-17977.
601.0000000000,-105.73,-13.012,-11.373,-15387.,-17977.
602.0000000000,-105.70,-13.009,-11.370,-15387.,-17977.
603.0000000000,-105.68,-13.007,-11.368,-15387.,-17977.
604.0000000000,-105.66,-13.006,-11.367,-15387.,-17977.
605.0000000000,-105.65,-13.005,-11.367,-15387.,-17977.
606.0000000000,-105.63,-13.004,-11.365,-15387.,-17976.
607.0000000000,-105.66,-13.008,-11.369,-15387.,-17976.
608.0000000000,-105.64,-13.007,-11.368,-15387.,-17976.
609.0000000000,-105.61,-13.005,-11.365,-15387.,-17976.
610.0000000000,-105.60,-13.003,-11.364,-15387.,-17976.
611.0000000000,-105.58,-13.001,-11.362,-15387.,-17976.
612.0000000000,-105.58,-13.001,-11.362,-15387.,-17976.
613.0000000000,-105.82,-13.030,-11.390,-15387.,-17976.
614.0000000000,-105.77,-13.027,-11.388,-15387.,-17976.
615.0000000000,-105.69,-13.017,-11.377,-15387.,-17976.
616.0000000000,-105.85,-13.033,-11.393,-15387.,-17976.
617.0000000000,-105.74,-13.021,-11.381,-15387.,-17976.
618.0000000000,-105.69,-13.013,-11.374,-15387.,-17976.
619.0000000000,-105.66,-13.008,-11.369,-15387.,-17976.
620.0000000000,-105.64,-13.005,-11.366,-15387.,-17976.
621.0000000000,-105.69,-13.011,-11.373,-15387.,-17975.
622.0000000000,-105.69,-13.014,-11.375,-15387.,-17975.
623.0000000000,-105.65,-13.008,-11.370,-15387.,-17975.
624.0000000000,-105.61,-13.004,-11.366,-15387.,-17975.
625.0000000000,-105.64,-13.007,-11.368,-15387.,-17975.
626.0000000000,-105.60,-13.003,-11.365,-15387.,-17975.
627.0000000000,-106.04,-13.053,-11.414,-15387.,-17975.
628.0000000000,-105.86,-13.037,-11.399,-15387.,-17975.
629.0000000000,-105.99,-13.049,-11.410,-15387.,-17975.
630.0000000000,-105.97,-13.046,-11.408,-15387.,-17975.
631.0000000000,-105.84,-13.029,-11.391,-15387.,-17975.
632.0000000000,-105.78,-13.018,-11.381,-15387.,-17975.
633.0000000000,-105.74,-13.012,-11.375,-15387.,-17975.
634.0000000000,-105.71,-13.009,-11.373,-15387.,-17975.
635.0000000000,-106.67,-13.119,-11.483,-15387.,-17975.
636.0000000000,-106.38,-13.096,-11.462,-15387.,-17975.
637.0000000000,-106.15,-13.063,-11.427,-15387.,-17975.
638.0000000000,-106.04,-13.041,-11.406,-15387.,-17975.
639.0000000000,-105.96,-13.028,-11.395,-15387.,-17975.
640.0000000000,-105.90,-13.019,-11.387,-15387.,-17974.
641.0000000000,-105.85,-13.014,-11.382,-15387.,-17974.
642.0000000000,-105.81,-13.010,-11.379,-15386.,-17974.
643.0000000000,-105.78,-13.007,-11.377,-15386.,-17974.
644.0000000000,-105.76,-13.005,-11.375,-15386.,-17974.
645.0000000000,-105.73,-13.003,-11.373,-15386.,-17974.
646.0000000000,-105.71,-13.002,-11.372,-15386.,-17974.
647.0000000000,-105.69,-13.001,-11.371,-15386.,-17974.
648.0000000000,-105.68,-12.999,-11.370,-15386.,-17973.
649.0000000000,-106.08,-13.046,-11.416,-15386.,-17973.
650.0000000000,-105.88,-13.029,-11.399,-15386.,-17973.
651.0000000000,-105.82,-13.018,-11.387,-15386.,-17973.
652.0000000000,-105.77,-13.011,-11.380,-15386.,-17973.
653.0000000000,-105.74,-13.006,-11.376,-15386.,-17973.
654.0000000000,-105.72,-13.003,-11.373,-15386.,-17973.
655.0000000000,-105.70,-13.001,-11.371,-15386.,-17973.
656.0000000000,-105.68,-12.999,-11.370,-15386.,-17973.
657.0000000000,-105.66,-12.998,-11.368,-15386.,-17973.
658.0000000000,-105.65,-12.997,-11.367,-15386.,-17972.
659.0000000000,-105.65,-12.998,-11.368,-15386.,-17972.
660.0000000000,-105.71,-13.006,-11.376,-15386.,-17972.
661.0000000000,-105.90,-13.029,-11.398,-15386.,-17972.
662.0000000000,-105.77,-13.016,-11.386,-15386.,-17972.
663.0000000000,-105.72,-13.008,-11.378,-15386.,-17972.
664.0000000000,-105.69,-13.003,-11.373,-15386.,-17972.
665.0000000000,-105.67,-12.999,-11.370,-15386.,-17972.
666.0000000000,-105.64,-12.997,-11.367,-15386.,-17972.
667.0000000000,-105.63,-12.995,-11.366,-15385.,-17972.
668.0000000000,-105.61,-12.993,-11.364,-15385.,-17972.
669.0000000000,-105.60,-12.992,-11.363,-15385.,-17971.
670.0000000000,-105.58,-12.991,-11.362,-15385.,-17971.
671.0000000000,-105.57,-12.990,-11.361,-15385.,-17971.
672.0000000000,-105.56,-12.990,-11.360,-15385.,-17971.
673.0000000000,-105.55,-12.989,-11.359,-15385.,-17971.
674.0000000000,-106.92,-13.146,-11.517,-15385.,-17971.
675.0000000000,-107.07,-13.177,-11.549,-15386.,-17972.
676.0000000000,-106.56,-13.116,-11.485,-15386.,-17972.
677.0000000000,-106.35,-13.077,-11.446,-15386.,-17972.
678.0000000000,-106.21,-13.050,-11.421,-15386.,-17972.
679.0000000000,-106.11,-13.033,-11.407,-15386.,-17972.
680.0000000000,-106.04,-13.022,-11.398,-15386.,-17972.
681.0000000000,-105.98,-13.015,-11.392,-15385.,-17971.
682.0000000000,-105.93,-13.010,-11.387,-15385.,-17971.
683.0000000000,-105.89,-13.006,-11.384,-15385.,-17971.
684.0000000000,-105.86,-13.004,-11.382,-15385.,-17971.
685.0000000000,-105.83,-13.002,-11.380,-15385.,-17971.
686.0000000000,-105.80,-13.000,-11.379,-15385.,-17971.
687.0000000000,-105.78,-12.999,-11.377,-15385.,-17970.
688.0000000000,-105.76,-12.997,-11.376,-15385.,-17970.
689.0000000000,-105.75,-12.996,-11.375,-15385.,-17970.
690.0000000000,-105.73,-12.995,-11.374,-15385.,-17970.
691.0000000000,-105.72,-12.995,-11.373,-15385.,-17970.
692.0000000000,-105.83,-13.009,-11.387,-15385.,-17970.
693.0000000000,-105.76,-13.003,-11.381,-15385.,-17970.
694.0000000000,-105.74,-12.999,-11.377,-15385.,-17970.
695.0000000000,-105.72,-12.996,-11.374,-15385.,-17970.
696.0000000000,-105.70,-12.994,-11.372,-15384.,-17969.
697.0000000000,-105.69,-12.993,-11.371,-15384.,-17969.
698.0000000000,-105.67,-12.992,-11.369,-15384.,-17969.
699.0000000000,-105.66,-12.991,-11.368,-15384.,-17969.
700.0000000000,-105.65,-12.990,-11.367,-15384.,-17969.
701.0000000000,-105.64,-12.989,-11.366,-15384.,-17969.
702.0000000000,-105.63,-12.988,-11.366,-15384.,-17969.
703.0000000000,-105.62,-12.987,-11.365,-15384.,-17969.
704.0000000000,-105.61,-12.987,-11.364,-15384.,-17969.
705.0000000000,-105.60,-12.986,-11.363,-15384.,-17968.
706.0000000000,-105.59,-12.985,-11.362,-15384.,-17968.
707.0000000000,-105.58,-12.985,-11.361,-15384.,-17968.
708.0000000000,-105.57,-12.984,-11.361,-15384.,-17968.
709.0000000000,-105.56,-12.984,-11.360,-15384.,-17968.
710.0000000000,-105.56,-12.984,-11.360,-15384.,-17968.
711.0000000000,-105.55,-12.983,-11.359,-15384.,-17968.
712.0000000000,-105.54,-12.982,-11.358,-15384.,-17968.
713.0000000000,-105.53,-12.981,-11.357,-15384.,-17968.
714.0000000000,-105.52,-12.980,-11.356,-15384.,-17968.
715.0000000000,-105.51,-12.980,-11.355,-15384.,-17968.
716.0000000000,-105.50,-12.979,-11.354,-15384.,-17967.
717.0000000000,-105.49,-12.978,-11.354,-15383.,-17967.
718.0000000000,-105.50,-12.980,-11.355,-15383.,-17967.
719.0000000000,-105.48,-12.979,-11.353,-15383.,-17967.
720.0000000000,-105.47,-12.977,-11.352,-15383.,-17967.
721.0000000000,-105.46,-12.976,-11.351,-15383.,-17967.
722.0000000000,-105.47,-12.978,-11.352,-15383.,-17967.
723.0000000000,-105.47,-12.979,-11.353,-15383.,-17967.
724.0000000000,-105.45,-12.977,-11.351,-15383.,-17967.
725.0000000000,-105.44,-12.975,-11.349,-15383.,-17967.
726.0000000000,-105.43,-12.974,-11.348,-15383.,-17967.
727.0000000000,-105.96,-13.035,-11.408,-15383.,-17967.
728.0000000000,-105.74,-13.015,-11.390,-15383.,-17967.
729.0000000000,-105.65,-13.001,-11.374,-15383.,-17967.
730.0000000000,-105.63,-12.995,-11.368,-15383.,-17967.
731.0000000000,-105.68,-13.000,-11.373,-15383.,-17967.
732.0000000000,-105.77,-13.010,-11.383,-15383.,-17967.
733.0000000000,-105.84,-13.018,-11.393,-15383.,-17967.
734.0000000000,-105.71,-13.002,-11.377,-15383.,-17966.
735.0000000000,-105.65,-12.992,-11.368,-15383.,-17966.
736.0000000000,-105.61,-12.986,-11.362,-15383.,-17966.
737.0000000000,-105.57,-12.981,-11.358,-15383.,-17966.
738.0000000000,-105.55,-12.978,-11.355,-15383.,-17966.
739.0000000000,-105.54,-12.978,-11.355,-15383.,-17966.
740.0000000000,-105.77,-13.006,-11.382,-15383.,-17966.
741.0000000000,-105.67,-12.997,-11.374,-15383.,-17966.
742.0000000000,-105.61,-12.988,-11.365,-15382.,-17965.
743.0000000000,-105.57,-12.982,-11.359,-15382.,-17965.
744.0000000000,-105.54,-12.978,-11.356,-15382.,-17965.
745.0000000000,-105.52,-12.975,-11.353,-15382.,-17965.
746.0000000000,-105.50,-12.973,-11.351,-15382.,-17965.
747.0000000000,-105.48,-12.972,-11.350,-15382.,-17965.
748.0000000000,-105.47,-12.970,-11.348,-15382.,-17965.
749.0000000000,-105.46,-12.969,-11.347,-15382.,-17964.
750.0000000000,-105.44,-12.968,-11.346,-15382.,-17964.
751.0000000000,-105.43,-12.968,-11.345,-15382.,-17964.
752.0000000000,-105.59,-12.987,-11.364,-15382.,-17964.
753.0000000000,-105.71,-13.003,-11.380,-15382.,-17964.
754.0000000000,-105.60,-12.991,-11.368,-15382.,-17964.
755.0000000000,-105.55,-12.983,-11.359,-15382.,-17964.
756.0000000000,-105.51,-12.977,-11.354,-15382.,-17964.
757.0000000000,-105.49,-12.973,-11.350,-15382.,-17964.
758.0000000000,-105.47,-12.970,-11.348,-15382.,-17964.
759.0000000000,-105.45,-12.968,-11.346,-15382.,-17964.
760.0000000000,-105.43,-12.966,-11.344,-15381.,-17963.
761.0000000000,-105.58,-12.984,-11.361,-15381.,-17963.
762.0000000000,-105.71,-13.002,-11.379,-15381.,-17963.
763.0000000000,-105.58,-12.988,-11.365,-15381.,-17963.
764.0000000000,-105.53,-12.979,-11.356,-15381.,-17963.
765.0000000000,-105.51,-12.975,-11.353,-15381.,-17963.
766.0000000000,-105.48,-12.971,-11.349,-15381.,-17963.
767.0000000000,-105.46,-12.968,-11.346,-15381.,-17963.
768.0000000000,-105.44,-12.965,-11.344,-15381.,-17963.
769.0000000000,-105.42,-12.964,-11.343,-15381.,-17963.
770.0000000000,-105.40,-12.962,-11.341,-15381.,-17962.
771.0000000000,-105.39,-12.961,-11.340,-15381.,-17962.
772.0000000000,-105.38,-12.960,-11.339,-15381.,-17962.
773.0000000000,-105.37,-12.959,-11.338,-15381.,-17962.
774.0000000000,-105.36,-12.959,-11.337,-15381.,-17962.
775.0000000000,-105.35,-12.958,-11.336,-15381.,-17962.
776.0000000000,-105.34,-12.957,-11.336,-15381.,-17962.
777.0000000000,-105.33,-12.957,-11.335,-15380.,-17962.
778.0000000000,-105.34,-12.959,-11.337,-15380.,-17961.
779.0000000000,-105.32,-12.957,-11.335,-15380.,-17961.
780.0000000000,-105.31,-12.956,-11.334,-15380.,-17961.
781.0000000000,-105.30,-12.955,-11.333,-15380.,-17961.
782.0000000000,-105.29,-12.954,-11.332,-15380.,-17961.
783.0000000000,-105.28,-12.953,-11.331,-15380.,-17961.
784.0000000000,-105.27,-12.952,-11.330,-15380.,-17961.
785.0000000000,-105.26,-12.952,-11.329,-15380.,-17961.
786.0000000000,-105.26,-12.951,-11.328,-15380.,-17961.
787.0000000000,-105.25,-12.950,-11.328,-15380.,-17960.
788.0000000000,-105.24,-12.950,-11.327,-15380.,-17960.
789.0000000000,-105.30,-12.957,-11.334,-15380.,-17960.
790.0000000000,-105.28,-12.956,-11.333,-15380.,-17960.
791.0000000000,-105.26,-12.955,-11.331,-15380.,-17960.
792.0000000000,-105.24,-12.952,-11.328,-15380.,-17960.
793.0000000000,-105.23,-12.950,-11.326,-15380.,-17960.
794.0000000000,-105.46,-12.976,-11.352,-15379.,-17960.
795.0000000000,-105.34,-12.965,-11.342,-15379.,-17960.
796.0000000000,-105.30,-12.958,-11.334,-15379.,-17960.
797.0000000000,-105.35,-12.963,-11.339,-15379.,-17960.
798.0000000000,-105.32,-12.960,-11.335,-15379.,-17960.
799.0000000000,-105.31,-12.959,-11.335,-15379.,-17960.
800.0000000000,-105.27,-12.954,-11.330,-15379.,-17959.
801.0000000000,-105.25,-12.950,-11.327,-15379.,-17959.
802.0000000000,-105.23,-12.948,-11.325,-15379.,-17959.
803.0000000000,-105.22,-12.946,-11.323,-15379.,-17959.
804.0000000000,-105.21,-12.945,-11.322,-15379.,-17959.
805.0000000000,-105.19,-12.944,-11.321,-15379.,-17959.
806.0000000000,-105.18,-12.943,-11.320,-15379.,-17958.
807.0000000000,-105.22,-12.948,-11.325,-15379.,-17958.
808.0000000000,-105.20,-12.946,-11.323,-15379.,-17958.
809.0000000000,-105.44,-12.975,-11.351,-15379.,-17958.
810.0000000000,-106.28,-13.072,-11.449,-15379.,-17958.
811.0000000000,-106.36,-13.089,-11.466,-15379.,-17959.
812.0000000000,-105.95,-13.038,-11.414,-15379.,-17959.
813.0000000000,-105.79,-13.006,-11.383,-15379.,-17959.
814.0000000000,-105.68,-12.986,-11.365,-15379.,-17959.
815.0000000000,-105.64,-12.978,-11.358,-15379.,-17959.
816.0000000000,-105.57,-12.969,-11.350,-15378.,-17958.
817.0000000000,-105.51,-12.962,-11.344,-15378.,-17958.
818.0000000000,-105.47,-12.958,-11.341,-15378.,-17958.
819.0000000000,-105.44,-12.954,-11.338,-15378.,-17957.
820.0000000000,-105.41,-12.952,-11.336,-15378.,-17957.
821.0000000000,-105.39,-12.950,-11.334,-15378.,-17957.
822.0000000000,-105.36,-12.949,-11.333,-15378.,-17957.
823.0000000000,-105.35,-12.948,-11.332,-15378.,-17957.
824.0000000000,-105.33,-12.947,-11.330,-15378.,-17957.
825.0000000000,-105.32,-12.946,-11.329,-15378.,-17957.
826.0000000000,-105.35,-12.951,-11.334,-15377.,-17957.
827.0000000000,-105.32,-12.948,-11.331,-15377.,-17956.
828.0000000000,-105.31,-12.948,-11.331,-15377.,-17956.
829.0000000000,-105.41,-12.960,-11.342,-15377.,-17956.
830.0000000000,-105.34,-12.953,-11.336,-15377.,-17956.
831.0000000000,-105.32,-12.949,-11.332,-15377.,-17956.
832.0000000000,-105.38,-12.956,-11.338,-15377.,-17956.
833.0000000000,-105.75,-12.999,-11.382,-15377.,-17956.
834.0000000000,-105.54,-12.978,-11.362,-15377.,-17956.
835.0000000000,-105.46,-12.966,-11.348,-15377.,-17956.
836.0000000000,-105.64,-12.983,-11.365,-15377.,-17956.
837.0000000000,-105.56,-12.975,-11.358,-15377.,-17956.
838.0000000000,-105.81,-13.002,-11.385,-15377.,-17956.
839.0000000000,-105.63,-12.983,-11.366,-15377.,-17956.
840.0000000000,-105.55,-12.969,-11.353,-15377.,-17956.
841.0000000000,-105.49,-12.961,-11.345,-15377.,-17955.
842.0000000000,-105.45,-12.955,-11.340,-15377.,-17955.
843.0000000000,-105.42,-12.951,-11.337,-15376.,-17955.
844.0000000000,-105.64,-12.976,-11.362,-15376.,-17955.
845.0000000000,-105.51,-12.964,-11.350,-15376.,-17955.
846.0000000000,-105.46,-12.957,-11.343,-15376.,-17955.
847.0000000000,-105.83,-12.998,-11.384,-15376.,-17955.
848.0000000000,-105.62,-12.978,-11.365,-15376.,-17955.
849.0000000000,-105.55,-12.966,-11.352,-15376.,-17955.
850.0000000000,-105.50,-12.958,-11.345,-15376.,-17954.
851.0000000000,-105.46,-12.953,-11.340,-15376.,-17954.
852.0000000000,-105.43,-12.950,-11.337,-15376.,-17954.
853.0000000000,-105.41,-12.947,-11.335,-15376.,-17954.
854.0000000000,-105.39,-12.945,-11.333,-15375.,-17954.
855.0000000000,-105.37,-12.944,-11.332,-15375.,-17954.
856.0000000000,-105.35,-12.943,-11.331,-15375.,-17953.
857.0000000000,-105.35,-12.943,-11.331,-15375.,-17953.
858.0000000000,-105.33,-12.942,-11.329,-15375.,-17953.
859.0000000000,-105.32,-12.941,-11.328,-15375.,-17953.
860.0000000000,-105.30,-12.940,-11.327,-15375.,-17953.
861.0000000000,-106.54,-13.081,-11.468,-15375.,-17953.
862.0000000000,-106.90,-13.135,-11.524,-15375.,-17954.
863.0000000000,-106.99,-13.145,-11.531,-15375.,-17954.
864.0000000000,-106.73,-13.106,-11.491,-15376.,-17955.
865.0000000000,-106.52,-13.069,-11.455,-15376.,-17955.
866.0000000000,-106.80,-13.089,-11.479,-15376.,-17955.
867.0000000000,-107.35,-13.149,-11.542,-15376.,-17955.
868.0000000000,-106.77,-13.084,-11.479,-15376.,-17955.
869.0000000000,-106.53,-13.044,-11.439,-15376.,-17955.
870.0000000000,-106.37,-13.018,-11.416,-15376.,-17955.
871.0000000000,-106.66,-13.048,-11.448,-15375.,-17954.
872.0000000000,-106.47,-13.031,-11.433,-15375.,-17954.
873.0000000000,-106.33,-13.013,-11.416,-15375.,-17954.
874.0000000000,-106.47,-13.027,-11.430,-15375.,-17954.
875.0000000000,-106.30,-13.010,-11.415,-15375.,-17953.
876.0000000000,-106.30,-13.009,-11.414,-15375.,-17953.
877.0000000000,-106.19,-12.996,-11.402,-15375.,-17953.
878.0000000000,-106.12,-12.987,-11.394,-15374.,-17952.
879.0000000000,-107.12,-13.101,-11.508,-15374.,-17952.
880.0000000000,-106.63,-13.058,-11.466,-15374.,-17953.
881.0000000000,-107.26,-13.122,-11.528,-15374.,-17953.
882.0000000000,-106.80,-13.070,-11.479,-15374.,-17953.
883.0000000000,-106.61,-13.039,-11.447,-15374.,-17952.
884.0000000000,-106.50,-13.019,-11.429,-15374.,-17952.
885.0000000000,-106.41,-13.006,-11.418,-15374.,-17952.
886.0000000000,-106.34,-12.998,-11.410,-15374.,-17952.
887.0000000000,-106.28,-12.992,-11.406,-15374.,-17952.
888.0000000000,-106.24,-12.988,-11.402,-15374.,-17952.
889.0000000000,-106.20,-12.985,-11.399,-15374.,-17951.
890.0000000000,-106.17,-12.983,-11.397,-15373.,-17951.
891.0000000000,-106.14,-12.981,-11.395,-15373.,-17951.
892.0000000000,-106.12,-12.980,-11.394,-15373.,-17951.
893.0000000000,-106.09,-12.978,-11.392,-15373.,-17950.
894.0000000000,-106.16,-12.988,-11.401,-15373.,-17950.
895.0000000000,-106.80,-13.063,-11.475,-15373.,-17950.
896.0000000000,-106.54,-13.041,-11.454,-15373.,-17951.
897.0000000000,-106.72,-13.057,-11.468,-15373.,-17951.
898.0000000000,-106.64,-13.046,-11.457,-15373.,-17951.
899.0000000000,-106.50,-13.026,-11.437,-15373.,-17951.
900.0000000000,-106.41,-13.012,-11.424,-15373.,-17950.
901.0000000000,-106.67,-13.039,-11.452,-15373.,-17950.
902.0000000000,-106.51,-13.023,-11.437,-15373.,-17950.
903.0000000000,-106.41,-13.009,-11.423,-15372.,-17950.
904.0000000000,-106.43,-13.010,-11.424,-15372.,-17950.
905.0000000000,-106.35,-13.001,-11.416,-15372.,-17950.
906.0000000000,-106.30,-12.994,-11.410,-15372.,-17950.
907.0000000000,-106.26,-12.990,-11.406,-15372.,-17949.
908.0000000000,-106.64,-13.035,-11.450,-15372.,-17949.
909.0000000000,-106.81,-13.059,-11.474,-15372.,-17949.
910.0000000000,-106.58,-13.035,-11.450,-15372.,-17949.
911.0000000000,-106.48,-13.017,-11.432,-15372.,-17949.
912.0000000000,-106.51,-13.017,-11.432,-15372.,-17949.
913.0000000000,-106.41,-13.006,-11.422,-15372.,-17949.
914.0000000000,-106.36,-12.998,-11.415,-15372.,-17949.
915.0000000000,-106.32,-12.993,-11.410,-15371.,-17949.
916.0000000000,-106.28,-12.990,-11.407,-15371.,-17949.
917.0000000000,-106.26,-12.987,-11.404,-15371.,-17948.
918.0000000000,-106.23,-12.985,-11.403,-15371.,-17948.
919.0000000000,-106.63,-13.033,-11.449,-15371.,-17948.
920.0000000000,-106.43,-13.014,-11.431,-15371.,-17948.
921.0000000000,-106.35,-13.003,-11.418,-15371.,-17948.
922.0000000000,-106.31,-12.995,-11.411,-15371.,-17948.
923.0000000000,-106.27,-12.990,-11.407,-15371.,-17948.
924.0000000000,-106.24,-12.987,-11.403,-15371.,-17948.
925.0000000000,-106.22,-12.985,-11.401,-15371.,-17947.
926.0000000000,-106.20,-12.983,-11.399,-15370.,-17947.
927.0000000000,-106.18,-12.981,-11.397,-15370.,-17947.
928.0000000000,-106.16,-12.980,-11.396,-15370.,-17947.
929.0000000000,-106.14,-12.979,-11.395,-15370.,-17947.
930.0000000000,-106.13,-12.978,-11.393,-15370.,-17947.
931.0000000000,-106.11,-12.977,-11.392,-15370.,-17947.
932.0000000000,-106.10,-12.977,-11.391,-15370.,-17946.
933.0000000000,-106.09,-12.976,-11.390,-15370.,-17946.
934.0000000000,-106.08,-12.975,-11.389,-15370.,-17946.
935.0000000000,-106.06,-12.974,-11.388,-15370.,-17946.
936.0000000000,-106.05,-12.974,-11.387,-15369.,-17946.
937.0000000000,-106.04,-12.973,-11.386,-15369.,-17946.
938.0000000000,-106.03,-12.972,-11.385,-15369.,-17946.
939.0000000000,-106.02,-12.972,-11.384,-15369.,-17946.
940.0000000000,-106.01,-12.971,-11.383,-15369.,-17945.
941.0000000000,-106.00,-12.970,-11.382,-15369.,-17945.
942.0000000000,-105.99,-12.969,-11.381,-15369.,-17945.
943.0000000000,-106.10,-12.983,-11.393,-15369.,-17945.
944.0000000000,-106.15,-12.992,-11.401,-15369.,-17945.
945.0000000000,-106.08,-12.983,-11.393,-15369.,-17945.
946.0000000000,-106.04,-12.977,-11.387,-15369.,-17945.
947.0000000000,-106.02,-12.973,-11.383,-15369.,-17945.
948.0000000000,-106.00,-12.971,-11.381,-15369.,-17945.
949.0000000000,-105.98,-12.969,-11.379,-15369.,-17944.
950.0000000000,-105.97,-12.967,-11.377,-15368.,-17944.
951.0000000000,-105.95,-12.966,-11.376,-15368.,-17944.
952.0000000000,-105.94,-12.965,-11.374,-15368.,-17944.
953.0000000000,-105.93,-12.964,-11.373,-15368.,-17944.
954.0000000000,-105.92,-12.963,-11.372,-15368.,-17944.
955.0000000000,-106.02,-12.977,-11.385,-15368.,-17944.
956.0000000000,-106.05,-12.982,-11.389,-15368.,-17944.
957.0000000000,-106.16,-12.996,-11.402,-15368.,-17943.
958.0000000000,-106.31,-13.013,-11.420,-15368.,-17944.
959.0000000000,-106.15,-12.995,-11.402,-15368.,-17943.
960.0000000000,-106.09,-12.983,-11.390,-15368.,-17943.
961.0000000000,-106.04,-12.976,-11.383,-15368.,-17943.
962.0000000000,-106.37,-13.012,-11.419,-15368.,-17943.
963.0000000000,-106.34,-13.012,-11.420,-15368.,-17943.
964.0000000000,-106.20,-12.995,-11.402,-15368.,-17943.
965.0000000000,-106.13,-12.984,-11.391,-15368.,-17943.
966.0000000000,-106.09,-12.976,-11.385,-15367.,-17943.
967.0000000000,-106.05,-12.971,-11.380,-15367.,-17942.
968.0000000000,-106.09,-12.977,-11.385,-15367.,-17942.
969.0000000000,-106.12,-12.982,-11.390,-15367.,-17942.
970.0000000000,-106.05,-12.974,-11.383,-15367.,-17942.
971.0000000000,-106.02,-12.969,-11.378,-15367.,-17942.
972.0000000000,-105.99,-12.966,-11.375,-15367.,-17942.
973.0000000000,-106.02,-12.970,-11.378,-15367.,-17942.
974.0000000000,-105.98,-12.966,-11.374,-15367.,-17941.
975.0000000000,-105.96,-12.963,-11.372,-15367.,-17941.
976.0000000000,-105.94,-12.961,-11.370,-15366.,-17941.
977.0000000000,-105.92,-12.960,-11.368,-15366.,-17941.
978.0000000000,-105.91,-12.958,-11.367,-15366.,-17941.
979.0000000000,-105.89,-12.957,-11.365,-15366.,-17941.
980.0000000000,-105.88,-12.956,-11.364,-15366.,-17940.
981.0000000000,-105.87,-12.955,-11.363,-15366.,-17940.
982.0000000000,-105.86,-12.955,-11.362,-15366.,-17940.
983.0000000000,-106.05,-12.978,-11.385,-15366.,-17940.
984.0000000000,-105.95,-12.969,-11.376,-15366.,-17940.
985.0000000000,-106.04,-12.978,-11.383,-15366.,-17940.
986.0000000000,-105.96,-12.968,-11.375,-15366.,-17940.
987.0000000000,-105.92,-12.963,-11.369,-15366.,-17940.
988.0000000000,-105.90,-12.959,-11.365,-15366.,-17940.
989.0000000000,-105.88,-12.956,-11.362,-15365.,-17939.
990.0000000000,-105.86,-12.954,-11.360,-15365.,-17939.
991.0000000000,-105.84,-12.953,-11.359,-15365.,-17939.
992.0000000000,-105.83,-12.951,-11.357,-15365.,-17939.
993.0000000000,-105.82,-12.950,-11.356,-15365.,-17939.
994.0000000000,-105.80,-12.949,-11.355,-15365.,-17939.
995.0000000000,-105.79,-12.948,-11.354,-15365.,-17939.
996.0000000000,-105.78,-12.948,-11.353,-15365.,-17938.
997.0000000000,-105.77,-12.947,-11.352,-15365.,-17938.
998.0000000000,-105.76,-12.946,-11.351,-15365.,-17938.
999.0000000000,-105.75,-12.945,-11.350,-15365.,-17938.
1000.000000000,-105.83,-12.955,-11.359,-15364.,-17938.
1001.000000000,-105.78,-12.951,-11.355,-15364.,-17938.
1002.000000000,-105.76,-12.948,-11.351,-15364.,-17938.
1003.000000000,-105.74,-12.946,-11.349,-15364.,-17938.
1004.000000000,-105.73,-12.944,-11.348,-15364.,-17937.
1005.000000000,-105.72,-12.943,-11.346,-15364.,-17937.
1006.000000000,-105.71,-12.942,-11.345,-15364.,-17937.
1007.000000000,-105.70,-12.941,-11.344,-15364.,-17937.
1008.000000000,-105.69,-12.941,-11.343,-15364.,-17937.
1009.000000000,-105.68,-12.940,-11.342,-15364.,-17937.
1010.000000000,-105.67,-12.939,-11.341,-15364.,-17937.
1011.000000000,-105.66,-12.939,-11.340,-15363.,-17937.
1012.000000000,-106.62,-13.048,-11.449,-15364.,-17937.
1013.000000000,-106.33,-13.026,-11.428,-15364.,-17937.
1014.000000000,-106.13,-12.996,-11.396,-15364.,-17937.
1015.000000000,-106.03,-12.977,-11.377,-15364.,-17937.
1016.000000000,-105.96,-12.965,-11.366,-15363.,-17937.
1017.000000000,-105.91,-12.957,-11.359,-15363.,-17937.
1018.000000000,-105.87,-12.952,-11.355,-15363.,-17937.
1019.000000000,-105.84,-12.948,-11.352,-15363.,-17936.
1020.000000000,-105.81,-12.946,-11.349,-15363.,-17936.
1021.000000000,-105.79,-12.944,-11.347,-15363.,-17936.
1022.000000000,-105.77,-12.942,-11.346,-15363.,-17936.
1023.000000000,-105.75,-12.941,-11.344,-15362.,-17936.
1024.000000000,-105.74,-12.940,-11.343,-15362.,-17936.
1025.000000000,-105.78,-12.947,-11.349,-15362.,-17936.
1026.000000000,-105.85,-12.956,-11.358,-15362.,-17936.
1027.000000000,-107.78,-13.177,-11.579,-15362.,-17936.
1028.000000000,-107.74,-13.192,-11.597,-15363.,-17937.
1029.000000000,-107.06,-13.105,-11.507,-15363.,-17937.
1030.000000000,-106.79,-13.052,-11.453,-15363.,-17937.
1031.000000000,-106.61,-13.018,-11.422,-15363.,-17937.
1032.000000000,-106.49,-12.997,-11.404,-15363.,-17937.
1033.000000000,-106.47,-12.993,-11.402,-15362.,-17936.
1034.000000000,-107.52,-13.114,-11.525,-15363.,-17937.
1035.000000000,-106.93,-13.058,-11.472,-15363.,-17937.
1036.000000000,-106.72,-13.025,-11.436,-15363.,-17937.
1037.000000000,-106.59,-13.003,-11.416,-15362.,-17936.
1038.000000000,-106.50,-12.989,-11.404,-15362.,-17936.
1039.000000000,-106.43,-12.980,-11.396,-15362.,-17935.
1040.000000000,-106.37,-12.974,-11.391,-15362.,-17935.
1041.000000000,-106.37,-12.976,-11.393,-15362.,-17935.
1042.000000000,-106.35,-12.977,-11.393,-15361.,-17935.
1043.000000000,-106.29,-12.971,-11.388,-15361.,-17934.
1044.000000000,-106.26,-12.967,-11.384,-15361.,-17934.
1045.000000000,-106.23,-12.964,-11.381,-15361.,-17934.
1046.000000000,-106.20,-12.962,-11.379,-15361.,-17934.
1047.000000000,-106.18,-12.961,-11.378,-15361.,-17934.
1048.000000000,-106.18,-12.963,-11.379,-15361.,-17933.
1049.000000000,-106.24,-12.971,-11.387,-15361.,-17933.
1050.000000000,-106.20,-12.968,-11.383,-15361.,-17933.
1051.000000000,-106.19,-12.968,-11.382,-15360.,-17933.
1052.000000000,-106.16,-12.963,-11.378,-15360.,-17933.
1053.000000000,-106.14,-12.960,-11.375,-15360.,-17933.
1054.000000000,-106.12,-12.958,-11.373,-15360.,-17933.
1055.000000000,-106.10,-12.956,-11.371,-15360.,-17932.
1056.000000000,-106.09,-12.955,-11.370,-15360.,-17932.
1057.000000000,-106.07,-12.954,-11.368,-15360.,-17932.
1058.000000000,-106.06,-12.953,-11.367,-15360.,-17932.
1059.000000000,-106.05,-12.952,-11.366,-15360.,-17932.
1060.000000000,-106.07,-12.956,-11.369,-15360.,-17932.
1061.000000000,-106.22,-12.974,-11.387,-15360.,-17932.
1062.000000000,-106.85,-13.049,-11.461,-15360.,-17932.
1063.000000000,-106.53,-13.018,-11.430,-15360.,-17932.
1064.000000000,-106.39,-12.995,-11.406,-15360.,-17932.
1065.000000000,-106.32,-12.980,-11.392,-15360.,-17932.
1066.000000000,-106.26,-12.971,-11.384,-15359.,-17932.
1067.000000000,-106.22,-12.965,-11.378,-15359.,-17932.
1068.000000000,-106.18,-12.961,-11.375,-15359.,-17931.
1069.000000000,-106.15,-12.958,-11.372,-15359.,-17931.
1070.000000000,-106.13,-12.956,-11.370,-15359.,-17931.
1071.000000000,-106.11,-12.954,-11.368,-15359.,-17931.
1072.000000000,-106.09,-12.953,-11.366,-15359.,-17931.
1073.000000000,-106.07,-12.952,-11.365,-15359.,-17930.
1074.000000000,-106.06,-12.951,-11.364,-15358.,-17930.
1075.000000000,-106.04,-12.950,-11.363,-15358.,-17930.
1076.000000000,-106.03,-12.949,-11.361,-15358.,-17930.
1077.000000000,-106.87,-13.046,-11.458,-15358.,-17930.
1078.000000000,-106.48,-13.010,-11.423,-15358.,-17930.
1079.000000000,-106.35,-12.989,-11.400,-15358.,-17930.
1080.000000000,-106.28,-12.976,-11.387,-15358.,-17930.
1081.000000000,-106.23,-12.967,-11.379,-15358.,-17930.
1082.000000000,-106.19,-12.961,-11.374,-15358.,-17930.
1083.000000000,-106.16,-12.957,-11.370,-15358.,-17930.
1084.000000000,-106.13,-12.955,-11.367,-15358.,-17930.
1085.000000000,-106.11,-12.953,-11.365,-15358.,-17929.
1086.000000000,-106.09,-12.951,-11.364,-15358.,-17929.
1087.000000000,-106.07,-12.950,-11.362,-15357.,-17929.
1088.000000000,-106.05,-12.949,-11.361,-15357.,-17929.
1089.000000000,-106.04,-12.948,-11.360,-15357.,-17929.
1090.000000000,-106.02,-12.947,-11.359,-15357.,-17929.
1091.000000000,-106.73,-13.029,-11.440,-15357.,-17929.
1092.000000000,-106.55,-13.016,-11.428,-15357.,-17929.
1093.000000000,-106.38,-12.992,-11.402,-15357.,-17929.
1094.000000000,-106.29,-12.976,-11.387,-15357.,-17929.
1095.000000000,-106.24,-12.967,-11.377,-15357.,-17929.
1096.000000000,-106.19,-12.960,-11.372,-15357.,-17929.
1097.000000000,-106.17,-12.958,-11.369,-15357.,-17929.
1098.000000000,-106.27,-12.970,-11.381,-15357.,-17928.
1099.000000000,-106.18,-12.962,-11.374,-15357.,-17928.
1100.000000000,-106.15,-12.957,-11.368,-15356.,-17928.
1101.000000000,-106.12,-12.953,-11.365,-15356.,-17928.
1102.000000000,-106.09,-12.950,-11.362,-15356.,-17928.
1103.000000000,-106.07,-12.948,-11.360,-15356.,-17928.
1104.000000000,-106.05,-12.947,-11.358,-15356.,-17927.
1105.000000000,-106.04,-12.946,-11.357,-15356.,-17927.
1106.000000000,-106.02,-12.945,-11.356,-15356.,-17927.
1107.000000000,-106.01,-12.944,-11.355,-15356.,-17927.
1108.000000000,-106.00,-12.943,-11.353,-15356.,-17927.
1109.000000000,-105.99,-12.942,-11.352,-15356.,-17927.
1110.000000000,-105.98,-12.942,-11.351,-15356.,-17927.
1111.000000000,-105.96,-12.941,-11.350,-15355.,-17927.
1112.000000000,-105.95,-12.940,-11.349,-15355.,-17926.
1113.000000000,-105.94,-12.939,-11.348,-15355.,-17926.
1114.000000000,-105.93,-12.939,-11.347,-15355.,-17926.
1115.000000000,-105.92,-12.938,-11.346,-15355.,-17926.
1116.000000000,-105.91,-12.937,-11.345,-15355.,-17926.
1117.000000000,-105.90,-12.937,-11.344,-15355.,-17926.
1118.000000000,-105.90,-12.936,-11.343,-15355.,-17926.
1119.000000000,-105.89,-12.936,-11.342,-15355.,-17926.
1120.000000000,-105.88,-12.935,-11.342,-15355.,-17925.
1121.000000000,-105.87,-12.934,-11.341,-15355.,-17925.
1122.000000000,-106.30,-12.985,-11.390,-15354.,-17925.
1123.000000000,-106.10,-12.966,-11.372,-15354.,-17925.
1124.000000000,-106.03,-12.955,-11.359,-15354.,-17925.
1125.000000000,-105.99,-12.947,-11.352,-15354.,-17925.
1126.000000000,-105.96,-12.942,-11.348,-15354.,-17925.
1127.000000000,-105.93,-12.939,-11.344,-15354.,-17925.
1128.000000000,-105.91,-12.937,-11.342,-15354.,-17925.
1129.000000000,-105.90,-12.935,-11.340,-15354.,-17925.
1130.000000000,-105.88,-12.934,-11.339,-15354.,-17924.
1131.000000000,-105.87,-12.933,-11.338,-15354.,-17924.
1132.000000000,-105.85,-12.932,-11.336,-15354.,-17924.
1133.000000000,-105.84,-12.931,-11.335,-15354.,-17924.
1134.000000000,-105.83,-12.930,-11.334,-15353.,-17924.
1135.000000000,-105.82,-12.929,-11.333,-15353.,-17924.
1136.000000000,-105.81,-12.929,-11.332,-15353.,-17924.
1137.000000000,-105.80,-12.928,-11.331,-15353.,-17924.
1138.000000000,-105.79,-12.927,-11.330,-15353.,-17923.
1139.000000000,-105.78,-12.927,-11.329,-15353.,-17923.
1140.000000000,-105.77,-12.926,-11.328,-15353.,-17923.
1141.000000000,-105.76,-12.925,-11.327,-15353.,-17923.
1142.000000000,-105.75,-12.925,-11.327,-15353.,-17923.
1143.000000000,-105.74,-12.924,-11.326,-15353.,-17923.
1144.000000000,-105.73,-12.923,-11.325,-15353.,-17923.
1145.000000000,-105.72,-12.923,-11.324,-15352.,-17923.
1146.000000000,-105.72,-12.922,-11.323,-15352.,-17922.
1147.000000000,-105.71,-12.922,-11.322,-15352.,-17922.
1148.000000000,-105.87,-12.941,-11.340,-15352.,-17922.
1149.000000000,-106.25,-12.987,-11.386,-15352.,-17922.
1150.000000000,-106.02,-12.963,-11.363,-15352.,-17922.
1151.000000000,-105.93,-12.949,-11.347,-15352.,-17922.
1152.000000000,-105.88,-12.939,-11.338,-15352.,-17922.
1153.000000000,-105.85,-12.933,-11.333,-15352.,-17922.
1154.000000000,-105.82,-12.929,-11.329,-15352.,-17922.
1155.000000000,-105.79,-12.926,-11.326,-15352.,-17922.
1156.000000000,-105.77,-12.924,-11.324,-15352.,-17922.
1157.000000000,-105.75,-12.923,-11.323,-15352.,-17921.
1158.000000000,-105.74,-12.921,-11.321,-15352.,-17921.
1159.000000000,-105.72,-12.920,-11.320,-15351.,-17921.
1160.000000000,-105.71,-12.919,-11.319,-15351.,-17921.
1161.000000000,-105.70,-12.918,-11.318,-15351.,-17921.
1162.000000000,-105.69,-12.918,-11.317,-15351.,-17921.
1163.000000000,-106.45,-13.006,-11.405,-15351.,-17921.
1164.000000000,-106.59,-13.030,-11.430,-15351.,-17921.
1165.000000000,-107.00,-13.075,-11.473,-15351.,-17921.
1166.000000000,-107.27,-13.104,-11.502,-15351.,-17922.
1167.000000000,-107.21,-13.093,-11.491,-15352.,-17922.
1168.000000000,-106.81,-13.036,-11.436,-15352.,-17922.
1169.000000000,-106.61,-13.001,-11.402,-15352.,-17922.
1170.000000000,-106.48,-12.978,-11.382,-15351.,-17922.
1171.000000000,-106.38,-12.964,-11.370,-15351.,-17921.
1172.000000000,-106.32,-12.957,-11.364,-15351.,-17921.
1173.000000000,-106.25,-12.949,-11.358,-15351.,-17920.
1174.000000000,-106.56,-12.986,-11.395,-15351.,-17921.
1175.000000000,-106.36,-12.968,-11.378,-15351.,-17920.
1176.000000000,-106.27,-12.956,-11.366,-15351.,-17920.
1177.000000000,-106.22,-12.949,-11.358,-15351.,-17920.
1178.000000000,-106.18,-12.944,-11.354,-15350.,-17920.
1179.000000000,-106.19,-12.946,-11.356,-15350.,-17919.
1180.000000000,-106.14,-12.942,-11.352,-15350.,-17919.
1181.000000000,-106.11,-12.939,-11.349,-15350.,-17919.
1182.000000000,-106.08,-12.936,-11.346,-15350.,-17919.
1183.000000000,-106.06,-12.934,-11.345,-15350.,-17919.
1184.000000000,-106.04,-12.933,-11.343,-15350.,-17918.
1185.000000000,-106.03,-12.932,-11.342,-15350.,-17918.
1186.000000000,-106.01,-12.931,-11.340,-15349.,-17918.
1187.000000000,-106.00,-12.932,-11.340,-15349.,-17918.
1188.000000000,-105.99,-12.930,-11.339,-15349.,-17918.
1189.000000000,-105.97,-12.929,-11.338,-15349.,-17918.
1190.000000000,-105.96,-12.928,-11.337,-15349.,-17918.
1191.000000000,-105.95,-12.927,-11.335,-15349.,-17917.
1192.000000000,-105.94,-12.927,-11.334,-15349.,-17917.
1193.000000000,-105.93,-12.926,-11.333,-15349.,-17917.
1194.000000000,-105.92,-12.925,-11.332,-15349.,-17917.
1195.000000000,-105.91,-12.925,-11.331,-15349.,-17917.
1196.000000000,-105.90,-12.924,-11.330,-15349.,-17917.
1197.000000000,-105.90,-12.925,-11.331,-15348.,-17916.
1198.000000000,-105.89,-12.924,-11.330,-15348.,-17916.
1199.000000000,-106.20,-12.960,-11.365,-15348.,-17916.
1200.000000000,-106.04,-12.946,-11.351,-15348.,-17916.
1201.000000000,-105.99,-12.937,-11.342,-15348.,-17916.
1202.000000000,-105.96,-12.932,-11.336,-15348.,-17916.
1203.000000000,-108.05,-13.170,-11.575,-15348.,-17917.
1204.000000000,-107.56,-13.135,-11.543,-15349.,-17917.
1205.000000000,-107.06,-13.066,-11.468,-15349.,-17917.
1206.000000000,-106.84,-13.022,-11.425,-15349.,-17917.
1207.000000000,-106.69,-12.993,-11.399,-15349.,-17917.
1208.000000000,-106.58,-12.975,-11.384,-15348.,-17917.
1209.000000000,-106.49,-12.963,-11.374,-15348.,-17917.
1210.000000000,-106.45,-12.959,-11.371,-15348.,-17916.
1211.000000000,-106.38,-12.952,-11.365,-15348.,-17916.
1212.000000000,-106.33,-12.947,-11.361,-15348.,-17916.
1213.000000000,-106.50,-12.968,-11.382,-15348.,-17916.
1214.000000000,-106.37,-12.957,-11.371,-15348.,-17916.
1215.000000000,-106.32,-12.950,-11.363,-15348.,-17915.
1216.000000000,-106.28,-12.945,-11.359,-15347.,-17915.
1217.000000000,-106.25,-12.942,-11.356,-15347.,-17915.
1218.000000000,-106.23,-12.941,-11.354,-15347.,-17915.
1219.000000000,-106.20,-12.938,-11.352,-15347.,-17915.
1220.000000000,-106.18,-12.937,-11.350,-15347.,-17914.
1221.000000000,-106.16,-12.935,-11.349,-15347.,-17914.
1222.000000000,-106.14,-12.934,-11.347,-15347.,-17914.
1223.000000000,-106.13,-12.933,-11.346,-15347.,-17914.
1224.000000000,-106.11,-12.932,-11.345,-15347.,-17914.
1225.000000000,-106.17,-12.940,-11.352,-15346.,-17914.
1226.000000000,-106.13,-12.936,-11.348,-15346.,-17914.
1227.000000000,-106.11,-12.934,-11.345,-15346.,-17914.
1228.000000000,-106.09,-12.932,-11.343,-15346.,-17913.
1229.000000000,-106.09,-12.932,-11.342,-15346.,-17913.
1230.000000000,-106.07,-12.931,-11.341,-15346.,-17913.
1231.000000000,-106.17,-12.943,-11.352,-15346.,-17913.
1232.000000000,-106.17,-12.945,-11.355,-15346.,-17913.
1233.000000000,-106.12,-12.939,-11.348,-15346.,-17913.
1234.000000000,-106.35,-12.965,-11.373,-15346.,-17913.
1235.000000000,-106.89,-13.028,-11.437,-15346.,-17913.
1236.000000000,-106.67,-13.008,-11.417,-15346.,-17913.
1237.000000000,-106.49,-12.981,-11.389,-15346.,-17913.
1238.000000000,-106.40,-12.963,-11.372,-15346.,-17913.
1239.000000000,-106.33,-12.952,-11.362,-15346.,-17913.
1240.000000000,-106.28,-12.945,-11.355,-15345.,-17913.
1241.000000000,-106.24,-12.940,-11.351,-15345.,-17913.
1242.000000000,-106.21,-12.937,-11.348,-15345.,-17913.
1243.000000000,-106.19,-12.935,-11.346,-15345.,-17912.
1244.000000000,-106.16,-12.933,-11.344,-15345.,-17912.
1245.000000000,-106.14,-12.931,-11.342,-15345.,-17912.
1246.000000000,-106.15,-12.934,-11.345,-15345.,-17912.
1247.000000000,-106.12,-12.932,-11.342,-15345.,-17912.
1248.000000000,-106.18,-12.939,-11.349,-15345.,-17912.
1249.000000000,-107.50,-13.092,-11.502,-15345.,-17912.
1250.000000000,-107.17,-13.068,-11.479,-15345.,-17912.
1251.000000000,-106.86,-13.024,-11.432,-15345.,-17912.
1252.000000000,-106.70,-12.993,-11.401,-15345.,-17912.
1253.000000000,-106.59,-12.973,-11.384,-15345.,-17912.
1254.000000000,-106.51,-12.961,-11.373,-15345.,-17912.
1255.000000000,-106.45,-12.952,-11.366,-15344.,-17912.
1256.000000000,-106.40,-12.947,-11.361,-15344.,-17912.
1257.000000000,-106.36,-12.943,-11.357,-15344.,-17911.
1258.000000000,-106.32,-12.940,-11.355,-15344.,-17911.
1259.000000000,-106.30,-12.938,-11.353,-15344.,-17911.
1260.000000000,-106.29,-12.939,-11.353,-15344.,-17911.
1261.000000000,-106.26,-12.937,-11.351,-15344.,-17911.
1262.000000000,-106.24,-12.935,-11.349,-15344.,-17911.
1263.000000000,-106.22,-12.934,-11.347,-15343.,-17910.
1264.000000000,-106.20,-12.932,-11.346,-15343.,-17910.
1265.000000000,-106.19,-12.932,-11.345,-15343.,-17910.
1266.000000000,-106.17,-12.931,-11.343,-15343.,-17910.
1267.000000000,-106.47,-12.966,-11.377,-15343.,-17910.
1268.000000000,-106.32,-12.952,-11.364,-15343.,-17910.
1269.000000000,-106.27,-12.944,-11.355,-15343.,-17910.
1270.000000000,-106.23,-12.939,-11.350,-15343.,-17910.
1271.000000000,-106.21,-12.935,-11.346,-15343.,-17910.
1272.000000000,-106.19,-12.932,-11.344,-15343.,-17909.
1273.000000000,-106.46,-12.965,-11.376,-15343.,-17909.
1274.000000000,-108.61,-13.214,-11.626,-15343.,-17910.
1275.000000000,-107.62,-13.123,-11.536,-15343.,-17910.
1276.000000000,-107.27,-13.062,-11.470,-15343.,-17911.
1277.000000000,-107.06,-13.020,-11.430,-15343.,-17911.
1278.000000000,-106.92,-12.994,-11.407,-15343.,-17911.
1279.000000000,-106.81,-12.977,-11.393,-15343.,-17910.
1280.000000000,-106.72,-12.966,-11.384,-15343.,-17910.
1281.000000000,-106.66,-12.959,-11.377,-15343.,-17910.
1282.000000000,-106.60,-12.954,-11.373,-15342.,-17909.
1283.000000000,-106.56,-12.950,-11.370,-15342.,-17909.
1284.000000000,-106.52,-12.948,-11.367,-15342.,-17909.
1285.000000000,-106.49,-12.946,-11.365,-15342.,-17909.
1286.000000000,-106.46,-12.944,-11.363,-15342.,-17909.
1287.000000000,-106.44,-12.943,-11.362,-15342.,-17908.
1288.000000000,-106.42,-12.942,-11.360,-15341.,-17908.
1289.000000000,-106.40,-12.940,-11.359,-15341.,-17908.
1290.000000000,-106.38,-12.940,-11.358,-15341.,-17908.
1291.000000000,-106.37,-12.939,-11.357,-15341.,-17908.
1292.000000000,-106.35,-12.938,-11.355,-15341.,-17907.
1293.000000000,-106.34,-12.937,-11.354,-15341.,-17907.
1294.000000000,-106.33,-12.936,-11.353,-15341.,-17907.
1295.000000000,-106.31,-12.936,-11.352,-15341.,-17907.
1296.000000000,-106.30,-12.935,-11.351,-15341.,-17907.
1297.000000000,-106.29,-12.934,-11.350,-15341.,-17907.
1298.000000000,-106.28,-12.934,-11.349,-15341.,-17907.
1299.000000000,-106.27,-12.933,-11.348,-15340.,-17907.
1300.000000000,-106.26,-12.932,-11.347,-15340.,-17907.
1301.000000000,-106.25,-12.932,-11.346,-15340.,-17907.
1302.000000000,-106.24,-12.931,-11.345,-15340.,-17906.
1303.000000000,-106.23,-12.932,-11.345,-15340.,-17906.
1304.000000000,-106.46,-12.959,-11.371,-15340.,-17906.
1305.000000000,-106.37,-12.952,-11.363,-15340.,-17906.
1306.000000000,-106.32,-12.944,-11.355,-15340.,-17906.
1307.000000000,-106.29,-12.940,-11.351,-15340.,-17906.
1308.000000000,-106.27,-12.936,-11.347,-15340.,-17906.
1309.000000000,-106.25,-12.933,-11.344,-15340.,-17906.
1310.000000000,-106.23,-12.931,-11.342,-15340.,-17906.
1311.000000000,-106.21,-12.930,-11.341,-15340.,-17906.
1312.000000000,-106.20,-12.928,-11.339,-15339.,-17906.
1313.000000000,-106.18,-12.927,-11.338,-15339.,-17905.
1314.000000000,-106.17,-12.927,-11.337,-15339.,-17905.
1315.000000000,-106.16,-12.926,-11.336,-15339.,-17905.
1316.000000000,-106.15,-12.925,-11.334,-15339.,-17905.
1317.000000000,-106.14,-12.924,-11.333,-15339.,-17905.
1318.000000000,-106.13,-12.924,-11.332,-15339.,-17905.
1319.000000000,-106.12,-12.923,-11.331,-15339.,-17905.
1320.000000000,-106.11,-12.922,-11.330,-15339.,-17905.
1321.000000000,-106.94,-13.019,-11.426,-15339.,-17905.
1322.000000000,-107.29,-13.068,-11.476,-15339.,-17905.
1323.000000000,-107.13,-13.049,-11.456,-15339.,-17905.
1324.000000000,-106.89,-13.014,-11.419,-15339.,-17906.
1325.000000000,-107.24,-13.044,-11.450,-15339.,-17906.
1326.000000000,-107.07,-13.024,-11.432,-15339.,-17906.
1327.000000000,-106.92,-13.000,-11.409,-15339.,-17906.
1328.000000000,-108.55,-13.181,-11.592,-15339.,-17906.
1329.000000000,-107.90,-13.121,-11.535,-15339.,-17906.
1330.000000000,-107.83,-13.100,-11.511,-15339.,-17906.
1331.000000000,-107.89,-13.095,-11.509,-15339.,-17906.
1332.000000000,-107.51,-13.045,-11.462,-15339.,-17906.
1333.000000000,-107.38,-13.021,-11.439,-15339.,-17906.
1334.000000000,-107.22,-12.998,-11.419,-15339.,-17906.
1335.000000000,-107.11,-12.984,-11.407,-15339.,-17906.
1336.000000000,-107.05,-12.978,-11.402,-15339.,-17905.
1337.000000000,-107.10,-12.986,-11.410,-15338.,-17905.
1338.000000000,-107.04,-12.982,-11.407,-15338.,-17905.
1339.000000000,-107.07,-12.987,-11.412,-15338.,-17904.
1340.000000000,-107.03,-12.984,-11.409,-15338.,-17904.
1341.000000000,-107.01,-12.982,-11.407,-15338.,-17904.
1342.000000000,-107.19,-13.002,-11.427,-15338.,-17904.
1343.000000000,-107.03,-12.986,-11.412,-15338.,-17904.
1344.000000000,-106.95,-12.975,-11.400,-15337.,-17904.
1345.000000000,-106.90,-12.968,-11.394,-15337.,-17903.
1346.000000000,-106.86,-12.963,-11.389,-15337.,-17903.
1347.000000000,-106.83,-12.959,-11.386,-15337.,-17903.
1348.000000000,-106.80,-12.957,-11.383,-15337.,-17903.
1349.000000000,-106.77,-12.955,-11.381,-15337.,-17902.
1350.000000000,-106.84,-12.964,-11.390,-15337.,-17902.
1351.000000000,-106.78,-12.959,-11.385,-15337.,-17902.
1352.000000000,-106.99,-12.983,-11.408,-15336.,-17902.
1353.000000000,-106.88,-12.974,-11.399,-15336.,-17902.
1354.000000000,-106.93,-12.978,-11.402,-15336.,-17902.
1355.000000000,-106.84,-12.968,-11.392,-15336.,-17902.
1356.000000000,-106.80,-12.962,-11.385,-15336.,-17902.
1357.000000000,-106.77,-12.957,-11.381,-15336.,-17902.
1358.000000000,-106.74,-12.954,-11.378,-15336.,-17901.
1359.000000000,-106.72,-12.952,-11.376,-15336.,-17901.
1360.000000000,-106.70,-12.950,-11.374,-15336.,-17901.
1361.000000000,-106.68,-12.949,-11.372,-15336.,-17901.
1362.000000000,-106.66,-12.948,-11.371,-15336.,-17901.
1363.000000000,-106.65,-12.947,-11.370,-15336.,-17901.
1364.000000000,-107.75,-13.074,-11.496,-15336.,-17901.
1365.000000000,-109.77,-13.320,-11.744,-15336.,-17902.
1366.000000000,-108.78,-13.221,-11.645,-15336.,-17903.
1367.000000000,-108.22,-13.131,-11.550,-15336.,-17903.
1368.000000000,-107.94,-13.074,-11.495,-15336.,-17903.
1369.000000000,-107.74,-13.038,-11.464,-15336.,-17903.
1370.000000000,-107.60,-13.015,-11.445,-15336.,-17903.
1371.000000000,-107.48,-13.001,-11.433,-15336.,-17903.
1372.000000000,-107.39,-12.991,-11.425,-15336.,-17902.
1373.000000000,-107.32,-12.984,-11.419,-15336.,-17901.
1374.000000000,-107.26,-12.980,-11.415,-15335.,-17901.
1375.000000000,-107.21,-12.976,-11.411,-15335.,-17901.
1376.000000000,-107.17,-12.973,-11.409,-15335.,-17900.
1377.000000000,-107.14,-12.972,-11.407,-15335.,-17900.
1378.000000000,-107.11,-12.970,-11.405,-15335.,-17900.
1379.000000000,-107.08,-12.969,-11.403,-15335.,-17899.
1380.000000000,-107.06,-12.967,-11.402,-15335.,-17899.
1381.000000000,-107.04,-12.966,-11.400,-15334.,-17899.
1382.000000000,-107.02,-12.965,-11.399,-15334.,-17899.
1383.000000000,-107.00,-12.964,-11.397,-15334.,-17899.
1384.000000000,-106.98,-12.963,-11.396,-15334.,-17899.
1385.000000000,-106.97,-12.962,-11.395,-15334.,-17898.
1386.000000000,-106.95,-12.962,-11.393,-15334.,-17898.
1387.000000000,-106.94,-12.961,-11.392,-15334.,-17898.
1388.000000000,-106.93,-12.960,-11.391,-15334.,-17898.
1389.000000000,-106.91,-12.959,-11.390,-15334.,-17898.
1390.000000000,-106.91,-12.959,-11.389,-15334.,-17898.
1391.000000000,-106.89,-12.958,-11.388,-15334.,-17898.
1392.000000000,-106.88,-12.957,-11.386,-15333.,-17898.
1393.000000000,-106.87,-12.957,-11.385,-15333.,-17898.
1394.000000000,-106.86,-12.956,-11.384,-15333.,-17897.
1395.000000000,-106.84,-12.955,-11.383,-15333.,-17897.
1396.000000000,-106.83,-12.954,-11.382,-15333.,-17897.
1397.000000000,-106.82,-12.954,-11.381,-15333.,-17897.
1398.000000000,-106.81,-12.953,-11.379,-15333.,-17897.
1399.000000000,-106.80,-12.952,-11.378,-15333.,-17897.
1400.000000000,-106.79,-12.951,-11.377,-15333.,-17897.
1401.000000000,-106.78,-12.951,-11.376,-15333.,-17897.
1402.000000000,-106.76,-12.950,-11.375,-15333.,-17896.
1403.000000000,-106.75,-12.949,-11.374,-15333.,-17896.
1404.000000000,-107.23,-13.005,-11.429,-15332.,-17896.
1405.000000000,-107.03,-12.987,-11.411,-15332.,-17896.
1406.000000000,-106.95,-12.976,-11.397,-15332.,-17896.
1407.000000000,-106.96,-12.974,-11.396,-15332.,-17896.
1408.000000000,-106.90,-12.965,-11.388,-15332.,-17896.
1409.000000000,-106.86,-12.960,-11.382,-15332.,-17896.
1410.000000000,-107.57,-13.040,-11.463,-15332.,-17896.
1411.000000000,-107.24,-13.011,-11.434,-15332.,-17896.
1412.000000000,-107.11,-12.990,-11.411,-15332.,-17896.
1413.000000000,-107.04,-12.976,-11.398,-15332.,-17896.
1414.000000000,-106.98,-12.967,-11.390,-15332.,-17896.
1415.000000000,-106.94,-12.962,-11.385,-15332.,-17896.
1416.000000000,-106.91,-12.958,-11.382,-15332.,-17896.
1417.000000000,-106.88,-12.955,-11.379,-15332.,-17895.
1418.000000000,-106.85,-12.953,-11.377,-15332.,-17895.
1419.000000000,-106.83,-12.951,-11.375,-15331.,-17895.
1420.000000000,-106.81,-12.950,-11.373,-15331.,-17895.
1421.000000000,-106.79,-12.948,-11.372,-15331.,-17895.
1422.000000000,-106.78,-12.947,-11.370,-15331.,-17895.
1423.000000000,-106.76,-12.946,-11.369,-15331.,-17895.
1424.000000000,-106.75,-12.946,-11.368,-15331.,-17894.
1425.000000000,-106.73,-12.945,-11.367,-15331.,-17894.
1426.000000000,-106.79,-12.952,-11.373,-15331.,-17894.
1427.000000000,-106.75,-12.949,-11.370,-15331.,-17894.
1428.000000000,-106.73,-12.946,-11.367,-15331.,-17894.
1429.000000000,-106.71,-12.944,-11.365,-15331.,-17894.
1430.000000000,-106.70,-12.943,-11.363,-15330.,-17894.
1431.000000000,-106.68,-12.942,-11.361,-15330.,-17894.
1432.000000000,-106.67,-12.941,-11.360,-15330.,-17894.
1433.000000000,-106.94,-12.973,-11.391,-15330.,-17894.
1434.000000000,-107.28,-13.015,-11.434,-15330.,-17894.
1435.000000000,-108.62,-13.171,-11.589,-15330.,-17894.
1436.000000000,-107.98,-13.108,-11.527,-15331.,-17895.
1437.000000000,-107.64,-13.052,-11.469,-15331.,-17895.
1438.000000000,-107.46,-13.017,-11.435,-15331.,-17895.
1439.000000000,-107.34,-12.995,-11.416,-15331.,-17895.
1440.000000000,-107.24,-12.981,-11.404,-15330.,-17894.
1441.000000000,-107.17,-12.971,-11.396,-15330.,-17894.
1442.000000000,-107.11,-12.965,-11.390,-15330.,-17894.
1443.000000000,-107.10,-12.966,-11.391,-15330.,-17893.
1444.000000000,-107.04,-12.961,-11.386,-15330.,-17893.
1445.000000000,-107.01,-12.957,-11.383,-15330.,-17893.
1446.000000000,-106.98,-12.956,-11.381,-15330.,-17893.
1447.000000000,-106.95,-12.953,-11.379,-15329.,-17893.
1448.000000000,-106.93,-12.951,-11.377,-15329.,-17893.
1449.000000000,-106.91,-12.950,-11.375,-15329.,-17893.
1450.000000000,-106.89,-12.949,-11.374,-15329.,-17892.
1451.000000000,-106.87,-12.948,-11.372,-15329.,-17892.
1452.000000000,-106.89,-12.952,-11.375,-15329.,-17892.
1453.000000000,-106.86,-12.949,-11.373,-15329.,-17892.
1454.000000000,-106.91,-12.956,-11.378,-15329.,-17892.
1455.000000000,-106.86,-12.951,-11.374,-15329.,-17892.
1456.000000000,-106.84,-12.948,-11.371,-15328.,-17892.
1457.000000000,-106.82,-12.946,-11.368,-15328.,-17892.
1458.000000000,-106.81,-12.945,-11.366,-15328.,-17891.
1459.000000000,-106.79,-12.943,-11.365,-15328.,-17891.
1460.000000000,-106.80,-12.945,-11.366,-15328.,-17891.
1461.000000000,-106.78,-12.944,-11.364,-15328.,-17891.
1462.000000000,-106.76,-12.942,-11.362,-15328.,-17891.
1463.000000000,-106.79,-12.946,-11.366,-15328.,-17891.
1464.000000000,-106.76,-12.943,-11.363,-15328.,-17891.
1465.000000000,-106.74,-12.941,-11.360,-15328.,-17891.
1466.000000000,-106.73,-12.940,-11.359,-15328.,-17891.
1467.000000000,-106.72,-12.939,-11.357,-15327.,-17890.
1468.000000000,-106.70,-12.938,-11.356,-15327.,-17890.
1469.000000000,-106.69,-12.937,-11.354,-15327.,-17890.
1470.000000000,-106.68,-12.936,-11.353,-15327.,-17890.
1471.000000000,-106.67,-12.935,-11.352,-15327.,-17890.
1472.000000000,-106.66,-12.934,-11.351,-15327.,-17890.
1473.000000000,-106.65,-12.934,-11.350,-15327.,-17890.
1474.000000000,-106.64,-12.933,-11.349,-15327.,-17890.
1475.000000000,-106.69,-12.940,-11.355,-15327.,-17890.
1476.000000000,-106.77,-12.951,-11.366,-15327.,-17890.
1477.000000000,-106.97,-12.975,-11.389,-15327.,-17890.
1478.000000000,-106.82,-12.959,-11.373,-15327.,-17890.
1479.000000000,-107.10,-12.989,-11.401,-15327.,-17890.
1480.000000000,-106.92,-12.968,-11.382,-15327.,-17890.
1481.000000000,-106.84,-12.956,-11.369,-15327.,-17890.
1482.000000000,-106.80,-12.948,-11.361,-15326.,-17890.
1483.000000000,-106.76,-12.942,-11.357,-15326.,-17890.
1484.000000000,-106.73,-12.939,-11.353,-15326.,-17889.
1485.000000000,-106.70,-12.936,-11.351,-15326.,-17889.
1486.000000000,-106.68,-12.934,-11.349,-15326.,-17889.
1487.000000000,-106.66,-12.933,-11.347,-15326.,-17889.
1488.000000000,-106.65,-12.931,-11.345,-15326.,-17889.
1489.000000000,-106.65,-12.933,-11.346,-15326.,-17889.
1490.000000000,-106.63,-12.932,-11.345,-15326.,-17889.
1491.000000000,-106.61,-12.930,-11.343,-15325.,-17888.
1492.000000000,-106.60,-12.929,-11.341,-15325.,-17888.
1493.000000000,-106.59,-12.928,-11.340,-15325.,-17888.
1494.000000000,-106.57,-12.927,-11.339,-15325.,-17888.
1495.000000000,-106.56,-12.926,-11.338,-15325.,-17888.
1496.000000000,-106.55,-12.925,-11.337,-15325.,-17888.
1497.000000000,-106.55,-12.927,-11.337,-15325.,-17888.
1498.000000000,-106.54,-12.925,-11.336,-15325.,-17888.
1499.000000000,-106.53,-12.924,-11.334,-15325.,-17888.
1500.000000000,-106.51,-12.923,-11.333,-15325.,-17888.
1501.000000000,-106.50,-12.923,-11.332,-15325.,-17887.
1502.000000000,-106.49,-12.922,-11.331,-15324.,-17887.
1503.000000000,-106.48,-12.921,-11.330,-15324.,-17887.
1504.000000000,-106.47,-12.920,-11.329,-15324.,-17887.
1505.000000000,-106.47,-12.920,-11.328,-15324.,-17887.
1506.000000000,-107.54,-13.044,-11.451,-15324.,-17887.
1507.000000000,-107.05,-12.999,-11.408,-15324.,-17887.
1508.000000000,-106.90,-12.972,-11.378,-15324.,-17888.
1509.000000000,-106.83,-12.958,-11.364,-15324.,-17888.
1510.000000000,-106.76,-12.946,-11.353,-15324.,-17887.
1511.000000000,-106.71,-12.938,-11.346,-15324.,-17887.
1512.000000000,-106.82,-12.951,-11.359,-15324.,-17887.
1513.000000000,-106.72,-12.941,-11.350,-15324.,-17887.
1514.000000000,-106.67,-12.935,-11.343,-15324.,-17887.
1515.000000000,-106.64,-12.930,-11.339,-15324.,-17887.
1516.000000000,-106.61,-12.928,-11.336,-15323.,-17886.
1517.000000000,-106.59,-12.925,-11.334,-15323.,-17886.
1518.000000000,-106.57,-12.924,-11.333,-15323.,-17886.
1519.000000000,-106.55,-12.922,-11.331,-15323.,-17886.
1520.000000000,-106.53,-12.921,-11.330,-15323.,-17886.
1521.000000000,-106.52,-12.920,-11.328,-15323.,-17886.
1522.000000000,-106.51,-12.920,-11.327,-15323.,-17886.
1523.000000000,-106.49,-12.919,-11.326,-15323.,-17885.
1524.000000000,-106.48,-12.918,-11.325,-15323.,-17885.
1525.000000000,-106.55,-12.927,-11.333,-15322.,-17885.
1526.000000000,-106.50,-12.923,-11.329,-15322.,-17885.
1527.000000000,-106.48,-12.920,-11.326,-15322.,-17885.
1528.000000000,-106.47,-12.918,-11.324,-15322.,-17885.
1529.000000000,-106.45,-12.917,-11.322,-15322.,-17885.
1530.000000000,-106.44,-12.916,-11.321,-15322.,-17885.
1531.000000000,-106.45,-12.918,-11.322,-15322.,-17885.
1532.000000000,-106.43,-12.916,-11.320,-15322.,-17885.
1533.000000000,-106.42,-12.914,-11.319,-15322.,-17885.
1534.000000000,-106.41,-12.914,-11.317,-15322.,-17885.
1535.000000000,-106.39,-12.913,-11.316,-15322.,-17884.
1536.000000000,-106.38,-12.912,-11.315,-15322.,-17884.
1537.000000000,-106.37,-12.911,-11.314,-15322.,-17884.
1538.000000000,-106.36,-12.910,-11.313,-15321.,-17884.
1539.000000000,-106.35,-12.910,-11.312,-15321.,-17884.
1540.000000000,-106.34,-12.909,-11.311,-15321.,-17884.
1541.000000000,-106.33,-12.908,-11.310,-15321.,-17884.
1542.000000000,-106.32,-12.908,-11.309,-15321.,-17884.
1543.000000000,-106.32,-12.907,-11.308,-15321.,-17883.
1544.000000000,-106.32,-12.909,-11.309,-15321.,-17883.
1545.000000000,-106.30,-12.907,-11.307,-15321.,-17883.
1546.000000000,-106.29,-12.906,-11.306,-15321.,-17883.
1547.000000000,-106.28,-12.905,-11.305,-15321.,-17883.
1548.000000000,-106.28,-12.904,-11.304,-15321.,-17883.
1549.000000000,-106.75,-12.960,-11.358,-15321.,-17883.
1550.000000000,-106.53,-12.939,-11.338,-15321.,-17883.
1551.000000000,-106.45,-12.927,-11.325,-15320.,-17883.
1552.000000000,-106.41,-12.919,-11.317,-15320.,-17883.
1553.000000000,-107.30,-13.019,-11.417,-15320.,-17883.
1554.000000000,-106.87,-12.978,-11.378,-15320.,-17883.
1555.000000000,-106.72,-12.953,-11.351,-15320.,-17883.
1556.000000000,-106.64,-12.937,-11.336,-15320.,-17883.
1557.000000000,-106.58,-12.927,-11.327,-15320.,-17883.
1558.000000000,-106.53,-12.921,-11.321,-15320.,-17882.
1559.000000000,-106.49,-12.916,-11.317,-15320.,-17882.
1560.000000000,-106.46,-12.913,-11.315,-15320.,-17882.
1561.000000000,-106.43,-12.911,-11.312,-15320.,-17882.
1562.000000000,-106.71,-12.944,-11.345,-15320.,-17882.
1563.000000000,-106.64,-12.941,-11.341,-15320.,-17882.
1564.000000000,-106.64,-12.940,-11.340,-15320.,-17881.
1565.000000000,-106.97,-12.976,-11.376,-15319.,-17882.
1566.000000000,-106.74,-12.952,-11.352,-15319.,-17882.
1567.000000000,-106.67,-12.940,-11.340,-15319.,-17881.
1568.000000000,-106.75,-12.946,-11.346,-15319.,-17881.
1569.000000000,-106.64,-12.933,-11.334,-15319.,-17881.
1570.000000000,-106.58,-12.925,-11.326,-15319.,-17881.
1571.000000000,-106.54,-12.919,-11.321,-15319.,-17881.
1572.000000000,-106.51,-12.915,-11.318,-15319.,-17881.
1573.000000000,-106.48,-12.913,-11.315,-15319.,-17880.
1574.000000000,-106.46,-12.911,-11.313,-15319.,-17880.
1575.000000000,-106.44,-12.909,-11.311,-15319.,-17880.
1576.000000000,-106.42,-12.908,-11.310,-15318.,-17880.
1577.000000000,-106.40,-12.907,-11.309,-15318.,-17880.
1578.000000000,-106.39,-12.906,-11.308,-15318.,-17880.
1579.000000000,-106.38,-12.905,-11.306,-15318.,-17880.
1580.000000000,-106.36,-12.904,-11.305,-15318.,-17879.
1581.000000000,-106.35,-12.904,-11.304,-15318.,-17879.
1582.000000000,-106.34,-12.903,-11.303,-15318.,-17879.
1583.000000000,-106.33,-12.902,-11.302,-15318.,-17879.
1584.000000000,-106.32,-12.902,-11.301,-15318.,-17879.
1585.000000000,-106.31,-12.901,-11.301,-15318.,-17879.
1586.000000000,-106.30,-12.900,-11.300,-15318.,-17879.
1587.000000000,-106.29,-12.900,-11.299,-15317.,-17879.
1588.000000000,-106.28,-12.899,-11.298,-15317.,-17879.
1589.000000000,-106.27,-12.899,-11.297,-15317.,-17878.
1590.000000000,-106.26,-12.898,-11.296,-15317.,-17878.
1591.000000000,-106.25,-12.897,-11.295,-15317.,-17878.
1592.000000000,-106.62,-12.941,-11.338,-15317.,-17878.
1593.000000000,-106.45,-12.925,-11.322,-15317.,-17878.
1594.000000000,-106.39,-12.915,-11.311,-15317.,-17878.
1595.000000000,-106.35,-12.908,-11.305,-15317.,-17878.
1596.000000000,-106.32,-12.904,-11.301,-15317.,-17878.
1597.000000000,-106.30,-12.901,-11.298,-15317.,-17878.
1598.000000000,-106.29,-12.901,-11.297,-15317.,-17877.
1599.000000000,-106.27,-12.899,-11.295,-15316.,-17877.
1600.000000000,-106.25,-12.897,-11.293,-15316.,-17877.
1601.000000000,-106.99,-12.982,-11.377,-15316.,-17877.
1602.000000000,-106.69,-12.957,-11.353,-15316.,-17877.
1603.000000000,-107.17,-13.007,-11.401,-15316.,-17877.
1604.000000000,-106.84,-12.969,-11.364,-15316.,-17878.
1605.000000000,-106.72,-12.948,-11.343,-15316.,-17878.
1606.000000000,-106.63,-12.932,-11.328,-15316.,-17877.
1607.000000000,-106.57,-12.921,-11.319,-15316.,-17877.
1608.000000000,-106.52,-12.914,-11.313,-15316.,-17877.
1609.000000000,-106.47,-12.910,-11.309,-15316.,-17877.
1610.000000000,-107.19,-12.993,-11.391,-15316.,-17877.
1611.000000000,-106.84,-12.962,-11.362,-15316.,-17877.
1612.000000000,-109.14,-13.220,-11.619,-15316.,-17877.
1613.000000000,-108.28,-13.141,-11.543,-15316.,-17878.
1614.000000000,-107.83,-13.070,-11.467,-15316.,-17878.
1615.000000000,-107.72,-13.037,-11.436,-15316.,-17878.
1616.000000000,-107.88,-13.046,-11.449,-15316.,-17878.
1617.000000000,-107.60,-13.011,-11.417,-15317.,-17878.
1618.000000000,-107.40,-12.982,-11.390,-15316.,-17878.
1619.000000000,-107.27,-12.964,-11.374,-15316.,-17878.
1620.000000000,-107.17,-12.952,-11.364,-15316.,-17877.
1621.000000000,-107.10,-12.943,-11.357,-15316.,-17877.
1622.000000000,-107.04,-12.938,-11.352,-15315.,-17876.
1623.000000000,-106.99,-12.934,-11.348,-15315.,-17876.
1624.000000000,-106.94,-12.931,-11.346,-15315.,-17876.
1625.000000000,-106.91,-12.929,-11.343,-15315.,-17875.
1626.000000000,-106.88,-12.927,-11.341,-15315.,-17875.
1627.000000000,-106.85,-12.926,-11.340,-15315.,-17875.
1628.000000000,-106.83,-12.925,-11.339,-15314.,-17875.
1629.000000000,-106.81,-12.924,-11.337,-15314.,-17875.
1630.000000000,-106.79,-12.923,-11.336,-15314.,-17874.
1631.000000000,-106.77,-12.922,-11.335,-15314.,-17874.
1632.000000000,-106.76,-12.921,-11.334,-15314.,-17874.
1633.000000000,-106.74,-12.920,-11.332,-15314.,-17874.
1634.000000000,-106.73,-12.919,-11.331,-15314.,-17874.
1635.000000000,-106.72,-12.919,-11.330,-15314.,-17874.
1636.000000000,-106.71,-12.920,-11.330,-15314.,-17874.
1637.000000000,-106.70,-12.919,-11.329,-15313.,-17874.
1638.000000000,-106.69,-12.918,-11.328,-15313.,-17873.
1639.000000000,-106.88,-12.941,-11.351,-15313.,-17873.
1640.000000000,-106.82,-12.937,-11.346,-15313.,-17873.
1641.000000000,-106.76,-12.929,-11.338,-15313.,-17873.
1642.000000000,-106.73,-12.924,-11.333,-15313.,-17873.
1643.000000000,-106.71,-12.921,-11.329,-15313.,-17873.
1644.000000000,-106.69,-12.919,-11.327,-15313.,-17873.
1645.000000000,-106.67,-12.917,-11.325,-15313.,-17873.
1646.000000000,-106.65,-12.915,-11.323,-15313.,-17873.
1647.000000000,-106.66,-12.918,-11.325,-15313.,-17873.
1648.000000000,-106.67,-12.920,-11.327,-15313.,-17873.
1649.000000000,-106.93,-12.951,-11.357,-15313.,-17872.
1650.000000000,-107.14,-12.978,-11.384,-15313.,-17873.
1651.000000000,-106.93,-12.955,-11.361,-15313.,-17873.
1652.000000000,-106.85,-12.940,-11.346,-15312.,-17873.
1653.000000000,-106.79,-12.931,-11.337,-15312.,-17872.
1654.000000000,-106.75,-12.925,-11.331,-15312.,-17872.
1655.000000000,-106.72,-12.921,-11.328,-15312.,-17872.
1656.000000000,-106.76,-12.926,-11.332,-15312.,-17872.
1657.000000000,-106.84,-12.937,-11.343,-15312.,-17872.
1658.000000000,-106.96,-12.952,-11.358,-15312.,-17872.
1659.000000000,-106.92,-12.949,-11.355,-15312.,-17872.
1660.000000000,-106.87,-12.942,-11.347,-15312.,-17872.
1661.000000000,-106.83,-12.937,-11.342,-15312.,-17872.
1662.000000000,-106.77,-12.928,-11.334,-15312.,-17871.
1663.000000000,-106.74,-12.923,-11.329,-15312.,-17871.
1664.000000000,-106.71,-12.919,-11.325,-15311.,-17871.
1665.000000000,-106.68,-12.917,-11.323,-15311.,-17871.
1666.000000000,-107.38,-12.997,-11.403,-15311.,-17871.
1667.000000000,-107.05,-12.967,-11.374,-15311.,-17871.
1668.000000000,-106.93,-12.948,-11.353,-15311.,-17871.
1669.000000000,-106.86,-12.936,-11.341,-15311.,-17871.
1670.000000000,-106.81,-12.928,-11.334,-15311.,-17871.
1671.000000000,-106.77,-12.923,-11.330,-15311.,-17870.
1672.000000000,-106.74,-12.919,-11.326,-15311.,-17870.
1673.000000000,-106.80,-12.927,-11.334,-15311.,-17870.
1674.000000000,-106.78,-12.927,-11.334,-15311.,-17870.
1675.000000000,-106.85,-12.936,-11.342,-15310.,-17870.
1676.000000000,-106.91,-12.944,-11.350,-15310.,-17870.
1677.000000000,-106.81,-12.932,-11.338,-15310.,-17870.
1678.000000000,-106.77,-12.927,-11.332,-15310.,-17870.
1679.000000000,-106.73,-12.921,-11.327,-15310.,-17869.
1680.000000000,-106.71,-12.918,-11.324,-15310.,-17869.
1681.000000000,-106.73,-12.921,-11.326,-15310.,-17869.
1682.000000000,-107.61,-13.022,-11.428,-15310.,-17869.
1683.000000000,-107.18,-12.982,-11.389,-15310.,-17869.
1684.000000000,-107.04,-12.960,-11.364,-15310.,-17870.
1685.000000000,-106.95,-12.943,-11.349,-15310.,-17869.
1686.000000000,-106.89,-12.933,-11.339,-15310.,-17869.
1687.000000000,-106.85,-12.926,-11.334,-15310.,-17869.
1688.000000000,-106.81,-12.922,-11.329,-15310.,-17869.
1689.000000000,-106.84,-12.927,-11.334,-15309.,-17868.
1690.000000000,-106.82,-12.926,-11.333,-15309.,-17868.
1691.000000000,-106.77,-12.921,-11.328,-15309.,-17868.
1692.000000000,-106.74,-12.918,-11.325,-15309.,-17868.
1693.000000000,-106.72,-12.915,-11.323,-15309.,-17868.
1694.000000000,-106.70,-12.913,-11.321,-15309.,-17868.
1695.000000000,-106.68,-12.912,-11.319,-15309.,-17868.
1696.000000000,-106.66,-12.911,-11.318,-15309.,-17867.
1697.000000000,-106.87,-12.936,-11.342,-15309.,-17867.
1698.000000000,-107.04,-12.958,-11.364,-15309.,-17867.
1699.000000000,-106.91,-12.945,-11.350,-15309.,-17867.
1700.000000000,-107.00,-12.953,-11.357,-15309.,-17867.
1701.000000000,-106.88,-12.938,-11.343,-15309.,-17867.
1702.000000000,-106.82,-12.928,-11.333,-15308.,-17867.
1703.000000000,-106.78,-12.921,-11.327,-15308.,-17867.
1704.000000000,-106.74,-12.917,-11.323,-15308.,-17867.
1705.000000000,-106.72,-12.914,-11.320,-15308.,-17867.
1706.000000000,-106.69,-12.912,-11.318,-15308.,-17866.
1707.000000000,-106.67,-12.910,-11.316,-15308.,-17866.
1708.000000000,-106.67,-12.911,-11.316,-15308.,-17866.
1709.000000000,-106.64,-12.909,-11.314,-15308.,-17866.
1710.000000000,-106.63,-12.908,-11.313,-15308.,-17866.
1711.000000000,-106.62,-12.907,-11.312,-15307.,-17866.
1712.000000000,-106.60,-12.906,-11.311,-15307.,-17865.
1713.000000000,-106.59,-12.905,-11.309,-15307.,-17865.
1714.000000000,-106.57,-12.904,-11.308,-15307.,-17865.
1715.000000000,-106.56,-12.903,-11.307,-15307.,-17865.
1716.000000000,-106.55,-12.902,-11.306,-15307.,-17865.
1717.000000000,-106.54,-12.901,-11.305,-15307.,-17865.
1718.000000000,-106.53,-12.901,-11.304,-15307.,-17865.
1719.000000000,-106.52,-12.900,-11.303,-15307.,-17864.
1720.000000000,-106.51,-12.899,-11.302,-15307.,-17864.
1721.000000000,-106.50,-12.899,-11.301,-15306.,-17864.
1722.000000000,-106.49,-12.898,-11.300,-15306.,-17864.
1723.000000000,-106.48,-12.897,-11.299,-15306.,-17864.
1724.000000000,-106.49,-12.899,-11.300,-15306.,-17864.
1725.000000000,-106.47,-12.898,-11.299,-15306.,-17864.
1726.000000000,-106.46,-12.897,-11.297,-15306.,-17864.
1727.000000000,-106.46,-12.898,-11.298,-15306.,-17864.
1728.000000000,-106.44,-12.896,-11.296,-15306.,-17864.
1729.000000000,-107.23,-12.987,-11.387,-15306.,-17864.
1730.000000000,-107.34,-13.008,-11.408,-15306.,-17864.
1731.000000000,-108.62,-13.153,-11.552,-15306.,-17864.
1732.000000000,-109.36,-13.244,-11.645,-15306.,-17865.
1733.000000000,-109.08,-13.207,-11.608,-15307.,-17866.
1734.000000000,-108.60,-13.132,-11.532,-15307.,-17866.
1735.000000000,-108.24,-13.069,-11.472,-15307.,-17866.
1736.000000000,-107.95,-13.021,-11.428,-15307.,-17866.
1737.000000000,-107.76,-12.990,-11.402,-15307.,-17866.
1738.000000000,-108.09,-13.025,-11.439,-15307.,-17866.
1739.000000000,-107.84,-13.002,-11.419,-15307.,-17866.
1740.000000000,-107.66,-12.978,-11.396,-15306.,-17865.
1741.000000000,-107.54,-12.963,-11.382,-15306.,-17865.
1742.000000000,-107.45,-12.953,-11.373,-15306.,-17864.
1743.000000000,-107.38,-12.946,-11.367,-15306.,-17864.
1744.000000000,-107.57,-12.970,-11.391,-15305.,-17863.
1745.000000000,-107.43,-12.958,-11.380,-15305.,-17863.
1746.000000000,-107.35,-12.949,-11.371,-15305.,-17863.
1747.000000000,-107.30,-12.943,-11.365,-15305.,-17863.
1748.000000000,-107.26,-12.938,-11.361,-15305.,-17862.
1749.000000000,-107.22,-12.935,-11.358,-15305.,-17862.
1750.000000000,-107.20,-12.934,-11.356,-15305.,-17862.
1751.000000000,-107.17,-12.932,-11.354,-15304.,-17862.
1752.000000000,-107.15,-12.930,-11.352,-15304.,-17862.
1753.000000000,-107.13,-12.929,-11.350,-15304.,-17861.
1754.000000000,-107.11,-12.928,-11.349,-15304.,-17861.
1755.000000000,-107.09,-12.927,-11.348,-15304.,-17861.
1756.000000000,-107.08,-12.926,-11.346,-15304.,-17861.
1757.000000000,-107.06,-12.925,-11.345,-15304.,-17861.
1758.000000000,-107.05,-12.924,-11.344,-15304.,-17861.
1759.000000000,-107.03,-12.924,-11.343,-15304.,-17861.
1760.000000000,-107.02,-12.923,-11.342,-15303.,-17860.
1761.000000000,-107.01,-12.922,-11.340,-15303.,-17860.
1762.000000000,-106.99,-12.921,-11.339,-15303.,-17860.
1763.000000000,-106.98,-12.921,-11.338,-15303.,-17860.
1764.000000000,-106.97,-12.920,-11.337,-15303.,-17860.
1765.000000000,-106.96,-12.919,-11.336,-15303.,-17860.
1766.000000000,-106.95,-12.919,-11.335,-15303.,-17860.
1767.000000000,-106.94,-12.918,-11.334,-15303.,-17860.
1768.000000000,-106.92,-12.918,-11.333,-15303.,-17860.
1769.000000000,-106.91,-12.917,-11.332,-15303.,-17860.
1770.000000000,-106.90,-12.916,-11.331,-15303.,-17859.
1771.000000000,-106.89,-12.916,-11.330,-15302.,-17859.
1772.000000000,-106.88,-12.915,-11.329,-15302.,-17859.
1773.000000000,-106.87,-12.914,-11.328,-15302.,-17859.
1774.000000000,-106.87,-12.915,-11.328,-15302.,-17859.
1775.000000000,-106.85,-12.914,-11.326,-15302.,-17859.
1776.000000000,-106.84,-12.913,-11.325,-15302.,-17859.
1777.000000000,-106.90,-12.921,-11.333,-15302.,-17859.
1778.000000000,-106.86,-12.917,-11.329,-15302.,-17859.
1779.000000000,-106.86,-12.918,-11.328,-15302.,-17859.
1780.000000000,-106.83,-12.915,-11.325,-15302.,-17859.
1781.000000000,-106.82,-12.913,-11.323,-15302.,-17858.
1782.000000000,-106.80,-12.911,-11.321,-15302.,-17858.
1783.000000000,-106.79,-12.910,-11.319,-15301.,-17858.
1784.000000000,-106.78,-12.909,-11.318,-15301.,-17858.
1785.000000000,-106.76,-12.908,-11.317,-15301.,-17858.
1786.000000000,-106.75,-12.907,-11.316,-15301.,-17858.
1787.000000000,-106.74,-12.906,-11.315,-15301.,-17858.
1788.000000000,-106.73,-12.905,-11.314,-15301.,-17858.
1789.000000000,-106.72,-12.905,-11.313,-15301.,-17858.
1790.000000000,-106.71,-12.904,-11.312,-15301.,-17858.
1791.000000000,-106.70,-12.903,-11.310,-15301.,-17857.
1792.000000000,-106.69,-12.903,-11.309,-15301.,-17857.
1793.000000000,-106.68,-12.902,-11.308,-15301.,-17857.
1794.000000000,-106.67,-12.901,-11.307,-15300.,-17857.
1795.000000000,-106.66,-12.901,-11.306,-15300.,-17857.
1796.000000000,-106.65,-12.900,-11.305,-15300.,-17857.
1797.000000000,-106.64,-12.899,-11.304,-15300.,-17857.
1798.000000000,-106.63,-12.899,-11.303,-15300.,-17857.
1799.000000000,-106.62,-12.898,-11.303,-15300.,-17857.
1800.000000000,-106.61,-12.897,-11.302,-15300.,-17856.
1801.000000000,-106.82,-12.922,-11.325,-15300.,-17856.
1802.000000000,-107.50,-13.003,-11.406,-15300.,-17857.
1803.000000000,-107.33,-12.991,-11.394,-15300.,-17857.
1804.000000000,-107.11,-12.959,-11.360,-15300.,-17857.
1805.000000000,-107.00,-12.938,-11.340,-15300.,-17857.
1806.000000000,-106.93,-12.925,-11.329,-15300.,-17857.
1807.000000000,-106.88,-12.917,-11.322,-15300.,-17856.
1808.000000000,-106.83,-12.912,-11.317,-15299.,-17856.
1809.000000000,-106.80,-12.908,-11.313,-15299.,-17856.
1810.000000000,-106.77,-12.905,-11.311,-15299.,-17856.
1811.000000000,-106.78,-12.907,-11.312,-15299.,-17856.
1812.000000000,-107.02,-12.937,-11.342,-15299.,-17856.
1813.000000000,-106.87,-12.923,-11.329,-15299.,-17855.
1814.000000000,-106.87,-12.922,-11.326,-15299.,-17855.
1815.000000000,-106.82,-12.914,-11.318,-15299.,-17855.
1816.000000000,-106.78,-12.908,-11.313,-15299.,-17855.
1817.000000000,-106.75,-12.905,-11.310,-15299.,-17855.
1818.000000000,-106.73,-12.904,-11.308,-15298.,-17855.
1819.000000000,-106.71,-12.901,-11.306,-15298.,-17855.
1820.000000000,-106.69,-12.899,-11.304,-15298.,-17855.
1821.000000000,-106.67,-12.898,-11.303,-15298.,-17854.
1822.000000000,-106.69,-12.901,-11.305,-15298.,-17854.
1823.000000000,-106.68,-12.901,-11.305,-15298.,-17854.
1824.000000000,-106.65,-12.899,-11.302,-15298.,-17854.
1825.000000000,-106.64,-12.897,-11.300,-15298.,-17854.
1826.000000000,-106.63,-12.895,-11.299,-15298.,-17854.
1827.000000000,-106.61,-12.894,-11.297,-15298.,-17854.
1828.000000000,-106.61,-12.895,-11.297,-15298.,-17854.
1829.000000000,-106.59,-12.893,-11.295,-15297.,-17853.
1830.000000000,-106.58,-12.892,-11.294,-15297.,-17853.
1831.000000000,-106.57,-12.891,-11.293,-15297.,-17853.
1832.000000000,-106.56,-12.890,-11.292,-15297.,-17853.
1833.000000000,-106.55,-12.889,-11.291,-15297.,-17853.
1834.000000000,-106.54,-12.888,-11.290,-15297.,-17853.
1835.000000000,-106.53,-12.888,-11.289,-15297.,-17853.
1836.000000000,-106.52,-12.887,-11.288,-15297.,-17853.
1837.000000000,-106.51,-12.886,-11.287,-15297.,-17853.
1838.000000000,-106.50,-12.886,-11.286,-15297.,-17853.
1839.000000000,-106.49,-12.885,-11.285,-15297.,-17852.
1840.000000000,-106.48,-12.884,-11.284,-15296.,-17852.
1841.000000000,-106.47,-12.884,-11.283,-15296.,-17852.
1842.000000000,-106.47,-12.886,-11.284,-15296.,-17852.
1843.000000000,-106.46,-12.884,-11.282,-15296.,-17852.
1844.000000000,-106.45,-12.883,-11.281,-15296.,-17852.
1845.000000000,-106.45,-12.884,-11.281,-15296.,-17852.
1846.000000000,-106.44,-12.884,-11.281,-15296.,-17852.
1847.000000000,-106.43,-12.883,-11.279,-15296.,-17852.
1848.000000000,-106.42,-12.881,-11.278,-15296.,-17851.
1849.000000000,-106.40,-12.880,-11.277,-15296.,-17851.
1850.000000000,-106.39,-12.879,-11.276,-15296.,-17851.
1851.000000000,-106.38,-12.878,-11.274,-15296.,-17851.
1852.000000000,-106.37,-12.877,-11.273,-15295.,-17851.
1853.000000000,-106.37,-12.877,-11.272,-15295.,-17851.
1854.000000000,-106.36,-12.876,-11.272,-15295.,-17851.
1855.000000000,-106.35,-12.875,-11.271,-15295.,-17850.
1856.000000000,-106.34,-12.875,-11.270,-15295.,-17850.
1857.000000000,-106.33,-12.874,-11.269,-15295.,-17850.
1858.000000000,-106.32,-12.873,-11.268,-15295.,-17850.
1859.000000000,-106.31,-12.873,-11.267,-15295.,-17850.
1860.000000000,-106.32,-12.875,-11.268,-15295.,-17850.
1861.000000000,-106.30,-12.873,-11.267,-15295.,-17850.
1862.000000000,-106.29,-12.872,-11.265,-15295.,-17850.
1863.000000000,-106.28,-12.871,-11.264,-15294.,-17850.
1864.000000000,-106.28,-12.872,-11.264,-15294.,-17849.
1865.000000000,-106.27,-12.871,-11.263,-15294.,-17849.
1866.000000000,-106.26,-12.870,-11.262,-15294.,-17849.
1867.000000000,-106.25,-12.869,-11.261,-15294.,-17849.
1868.000000000,-106.24,-12.868,-11.260,-15294.,-17849.
1869.000000000,-106.23,-12.867,-11.259,-15294.,-17849.
1870.000000000,-106.27,-12.873,-11.264,-15294.,-17849.
1871.000000000,-106.26,-12.873,-11.264,-15294.,-17849.
1872.000000000,-106.24,-12.870,-11.261,-15294.,-17849.
1873.000000000,-106.22,-12.868,-11.258,-15294.,-17848.
1874.000000000,-106.21,-12.866,-11.257,-15294.,-17848.
1875.000000000,-106.20,-12.865,-11.255,-15293.,-17848.
1876.000000000,-106.27,-12.874,-11.263,-15293.,-17848.
1877.000000000,-106.45,-12.897,-11.286,-15293.,-17848.
1878.000000000,-107.24,-12.989,-11.378,-15293.,-17848.
1879.000000000,-106.86,-12.952,-11.342,-15293.,-17849.
1880.000000000,-106.68,-12.923,-11.311,-15293.,-17849.
1881.000000000,-106.60,-12.907,-11.295,-15293.,-17849.
1882.000000000,-106.53,-12.894,-11.283,-15293.,-17848.
1883.000000000,-106.47,-12.885,-11.276,-15293.,-17848.
1884.000000000,-106.43,-12.879,-11.271,-15293.,-17848.
1885.000000000,-106.39,-12.876,-11.268,-15293.,-17848.
1886.000000000,-106.41,-12.879,-11.271,-15293.,-17848.
1887.000000000,-106.37,-12.875,-11.267,-15293.,-17847.
1888.000000000,-106.34,-12.872,-11.264,-15292.,-17847.
1889.000000000,-106.32,-12.870,-11.262,-15292.,-17847.
1890.000000000,-106.30,-12.868,-11.261,-15292.,-17847.
1891.000000000,-106.28,-12.867,-11.259,-15292.,-17847.
1892.000000000,-106.27,-12.866,-11.258,-15292.,-17847.
1893.000000000,-106.25,-12.865,-11.257,-15292.,-17847.
1894.000000000,-106.24,-12.864,-11.256,-15292.,-17846.
1895.000000000,-106.23,-12.863,-11.255,-15292.,-17846.
1896.000000000,-106.22,-12.863,-11.254,-15292.,-17846.
1897.000000000,-106.21,-12.862,-11.253,-15291.,-17846.
1898.000000000,-106.20,-12.861,-11.252,-15291.,-17846.
1899.000000000,-106.19,-12.861,-11.251,-15291.,-17846.
1900.000000000,-106.18,-12.860,-11.250,-15291.,-17846.
1901.000000000,-106.17,-12.860,-11.249,-15291.,-17846.
1902.000000000,-106.16,-12.859,-11.249,-15291.,-17846.
1903.000000000,-106.15,-12.858,-11.248,-15291.,-17845.
1904.000000000,-106.14,-12.858,-11.247,-15291.,-17845.
1905.000000000,-106.13,-12.857,-11.246,-15291.,-17845.
1906.000000000,-106.12,-12.857,-11.245,-15291.,-17845.
1907.000000000,-106.11,-12.856,-11.244,-15291.,-17845.
1908.000000000,-106.10,-12.856,-11.243,-15290.,-17845.
1909.000000000,-106.09,-12.855,-11.243,-15290.,-17845.
1910.000000000,-106.09,-12.854,-11.242,-15290.,-17845.
1911.000000000,-106.08,-12.854,-11.241,-15290.,-17845.
1912.000000000,-106.07,-12.853,-11.240,-15290.,-17844.
1913.000000000,-106.11,-12.859,-11.245,-15290.,-17844.
1914.000000000,-106.08,-12.856,-11.242,-15290.,-17844.
1915.000000000,-106.06,-12.854,-11.240,-15290.,-17844.
1916.000000000,-106.05,-12.853,-11.239,-15290.,-17844.
1917.000000000,-106.04,-12.852,-11.237,-15290.,-17844.
1918.000000000,-106.03,-12.851,-11.236,-15290.,-17844.
1919.000000000,-106.02,-12.850,-11.235,-15290.,-17844.
1920.000000000,-106.01,-12.849,-11.234,-15289.,-17844.
1921.000000000,-106.00,-12.849,-11.234,-15289.,-17843.
1922.000000000,-105.99,-12.848,-11.233,-15289.,-17843.
1923.000000000,-105.98,-12.848,-11.232,-15289.,-17843.
1924.000000000,-105.98,-12.847,-11.231,-15289.,-17843.
1925.000000000,-105.97,-12.846,-11.230,-15289.,-17843.
1926.000000000,-105.96,-12.846,-11.229,-15289.,-17843.
1927.000000000,-105.95,-12.845,-11.229,-15289.,-17843.
1928.000000000,-105.94,-12.845,-11.228,-15289.,-17843.
1929.000000000,-105.93,-12.844,-11.227,-15289.,-17842.
1930.000000000,-105.95,-12.847,-11.229,-15289.,-17842.
1931.000000000,-105.93,-12.845,-11.227,-15288.,-17842.
1932.000000000,-105.92,-12.844,-11.226,-15288.,-17842.
1933.000000000,-105.91,-12.843,-11.225,-15288.,-17842.
1934.000000000,-105.90,-12.842,-11.224,-15288.,-17842.
1935.000000000,-105.89,-12.841,-11.223,-15288.,-17842.
1936.000000000,-105.88,-12.841,-11.222,-15288.,-17842.
1937.000000000,-105.88,-12.840,-11.222,-15288.,-17842.
1938.000000000,-105.88,-12.842,-11.222,-15288.,-17841.
1939.000000000,-105.87,-12.841,-11.221,-15288.,-17841.
1940.000000000,-105.86,-12.840,-11.220,-15288.,-17841.
1941.000000000,-105.85,-12.839,-11.219,-15288.,-17841.
1942.000000000,-105.99,-12.856,-11.235,-15287.,-17841.
1943.000000000,-105.91,-12.849,-11.228,-15287.,-17841.
1944.000000000,-105.88,-12.844,-11.224,-15287.,-17841.
1945.000000000,-105.87,-12.841,-11.221,-15287.,-17841.
1946.000000000,-105.85,-12.839,-11.218,-15287.,-17841.
1947.000000000,-105.84,-12.838,-11.217,-15287.,-17841.
1948.000000000,-105.82,-12.837,-11.216,-15287.,-17840.
1949.000000000,-105.86,-12.842,-11.220,-15287.,-17840.
1950.000000000,-106.88,-12.959,-11.337,-15287.,-17840.
1951.000000000,-106.56,-12.934,-11.313,-15287.,-17841.
1952.000000000,-106.34,-12.900,-11.277,-15287.,-17841.
1953.000000000,-106.23,-12.879,-11.257,-15287.,-17841.
1954.000000000,-106.16,-12.865,-11.245,-15287.,-17841.
1955.000000000,-106.10,-12.857,-11.237,-15287.,-17840.
1956.000000000,-106.06,-12.851,-11.233,-15287.,-17840.
1957.000000000,-106.02,-12.847,-11.229,-15286.,-17840.
1958.000000000,-105.99,-12.845,-11.227,-15286.,-17840.
1959.000000000,-105.97,-12.843,-11.225,-15286.,-17839.
1960.000000000,-105.94,-12.841,-11.223,-15286.,-17839.
1961.000000000,-105.93,-12.840,-11.222,-15286.,-17839.
1962.000000000,-105.91,-12.839,-11.221,-15286.,-17839.
1963.000000000,-105.89,-12.838,-11.220,-15286.,-17839.
1964.000000000,-105.89,-12.839,-11.220,-15286.,-17839.
1965.000000000,-105.87,-12.837,-11.219,-15286.,-17839.
1966.000000000,-105.96,-12.848,-11.229,-15285.,-17838.
1967.000000000,-106.91,-12.958,-11.339,-15285.,-17839.
1968.000000000,-106.47,-12.917,-11.299,-15286.,-17839.
1969.000000000,-106.30,-12.890,-11.269,-15286.,-17839.
1970.000000000,-106.21,-12.872,-11.253,-15285.,-17839.
1971.000000000,-106.15,-12.861,-11.243,-15285.,-17839.
1972.000000000,-106.10,-12.854,-11.236,-15285.,-17838.
1973.000000000,-106.06,-12.849,-11.232,-15285.,-17838.
1974.000000000,-106.03,-12.846,-11.229,-15285.,-17838.
1975.000000000,-106.00,-12.843,-11.227,-15285.,-17838.
1976.000000000,-105.98,-12.842,-11.225,-15285.,-17838.
1977.000000000,-105.96,-12.840,-11.224,-15285.,-17837.
1978.000000000,-105.94,-12.839,-11.223,-15284.,-17837.
1979.000000000,-105.93,-12.838,-11.222,-15284.,-17837.
1980.000000000,-105.91,-12.837,-11.221,-15284.,-17837.
1981.000000000,-105.95,-12.843,-11.226,-15284.,-17837.
1982.000000000,-105.92,-12.840,-11.223,-15284.,-17837.
1983.000000000,-105.90,-12.838,-11.221,-15284.,-17837.
1984.000000000,-105.88,-12.837,-11.219,-15284.,-17837.
1985.000000000,-105.87,-12.835,-11.218,-15284.,-17836.
1986.000000000,-105.86,-12.834,-11.217,-15284.,-17836.
1987.000000000,-105.85,-12.834,-11.216,-15284.,-17836.
1988.000000000,-105.84,-12.833,-11.215,-15284.,-17836.
1989.000000000,-105.83,-12.832,-11.214,-15284.,-17836.
1990.000000000,-105.82,-12.832,-11.213,-15283.,-17836.
1991.000000000,-105.81,-12.831,-11.212,-15283.,-17836.
1992.000000000,-105.80,-12.830,-11.211,-15283.,-17836.
1993.000000000,-105.79,-12.830,-11.211,-15283.,-17836.
1994.000000000,-105.78,-12.829,-11.210,-15283.,-17835.
1995.000000000,-105.78,-12.829,-11.209,-15283.,-17835.
1996.000000000,-105.84,-12.837,-11.217,-15283.,-17835.
1997.000000000,-105.80,-12.834,-11.213,-15283.,-17835.
1998.000000000,-105.78,-12.831,-11.210,-15283.,-17835.
1999.000000000,-105.78,-12.832,-11.210,-15283.,-17835.
2000.000000000,-105.76,-12.830,-11.208,-15283.,-17835.
2001.000000000,-105.75,-12.828,-11.207,-15282.,-17835.
2002.000000000,-105.73,-12.827,-11.206,-15282.,-17834.
2003.000000000,-105.72,-12.826,-11.204,-15282.,-17834.
2004.000000000,-105.71,-12.825,-11.204,-15282.,-17834.
2005.000000000,-105.70,-12.825,-11.203,-15282.,-17834.
2006.000000000,-105.70,-12.824,-11.202,-15282.,-17834.
2007.000000000,-105.74,-12.831,-11.208,-15282.,-17834.
2008.000000000,-105.71,-12.827,-11.205,-15282.,-17834.
2009.000000000,-105.69,-12.825,-11.202,-15282.,-17834.
2010.000000000,-105.68,-12.824,-11.201,-15282.,-17833.
2011.000000000,-105.67,-12.823,-11.199,-15282.,-17833.
2012.000000000,-105.77,-12.835,-11.211,-15281.,-17833.
2013.000000000,-105.89,-12.851,-11.227,-15281.,-17833.
2014.000000000,-106.22,-12.890,-11.265,-15281.,-17833.
2015.000000000,-106.44,-12.917,-11.293,-15281.,-17833.
2016.000000000,-106.35,-12.906,-11.282,-15282.,-17834.
2017.000000000,-106.47,-12.915,-11.290,-15282.,-17834.
2018.000000000,-106.23,-12.883,-11.260,-15282.,-17834.
2019.000000000,-106.12,-12.864,-11.242,-15281.,-17833.
2020.000000000,-106.05,-12.852,-11.231,-15281.,-17833.
2021.000000000,-105.99,-12.844,-11.224,-15281.,-17833.
2022.000000000,-105.95,-12.839,-11.219,-15281.,-17833.
2023.000000000,-105.91,-12.835,-11.216,-15281.,-17832.
2024.000000000,-105.88,-12.832,-11.214,-15281.,-17832.
2025.000000000,-105.86,-12.830,-11.212,-15281.,-17832.
2026.000000000,-105.83,-12.829,-11.210,-15280.,-17832.
2027.000000000,-105.81,-12.827,-11.209,-15280.,-17832.
2028.000000000,-105.80,-12.826,-11.208,-15280.,-17831.
2029.000000000,-105.78,-12.826,-11.207,-15280.,-17831.
2030.000000000,-105.77,-12.825,-11.206,-15280.,-17831.
2031.000000000,-105.76,-12.824,-11.205,-15280.,-17831.
2032.000000000,-105.74,-12.823,-11.204,-15280.,-17831.
2033.000000000,-105.73,-12.823,-11.203,-15280.,-17831.
2034.000000000,-105.72,-12.822,-11.202,-15280.,-17831.
2035.000000000,-105.71,-12.821,-11.201,-15280.,-17831.
2036.000000000,-105.70,-12.821,-11.201,-15280.,-17831.
2037.000000000,-105.69,-12.820,-11.200,-15279.,-17830.
2038.000000000,-106.72,-12.938,-11.317,-15279.,-17831.
2039.000000000,-106.28,-12.899,-11.280,-15280.,-17831.
2040.000000000,-106.12,-12.873,-11.250,-15280.,-17831.
2041.000000000,-106.03,-12.856,-11.234,-15279.,-17831.
2042.000000000,-105.97,-12.845,-11.224,-15279.,-17831.
2043.000000000,-105.92,-12.838,-11.218,-15279.,-17830.
2044.000000000,-105.89,-12.833,-11.214,-15279.,-17830.
2045.000000000,-105.85,-12.830,-11.211,-15279.,-17830.
2046.000000000,-105.83,-12.828,-11.209,-15279.,-17830.
2047.000000000,-105.81,-12.826,-11.208,-15279.,-17830.
2048.000000000,-105.79,-12.825,-11.207,-15279.,-17829.
2049.000000000,-106.17,-12.869,-11.250,-15279.,-17829.
2050.000000000,-106.25,-12.884,-11.265,-15279.,-17829.
2051.000000000,-106.43,-12.904,-11.285,-15279.,-17829.
2052.000000000,-106.28,-12.886,-11.267,-15279.,-17829.
2053.000000000,-106.14,-12.865,-11.246,-15279.,-17829.
2054.000000000,-106.06,-12.852,-11.233,-15278.,-17829.
2055.000000000,-106.01,-12.843,-11.225,-15278.,-17829.
2056.000000000,-105.96,-12.837,-11.220,-15278.,-17829.
2057.000000000,-105.93,-12.833,-11.217,-15278.,-17829.
2058.000000000,-105.99,-12.841,-11.225,-15278.,-17828.
2059.000000000,-106.09,-12.855,-11.238,-15278.,-17828.
2060.000000000,-105.98,-12.844,-11.228,-15278.,-17828.
2061.000000000,-105.94,-12.837,-11.221,-15278.,-17828.
2062.000000000,-105.90,-12.833,-11.217,-15278.,-17828.
2063.000000000,-105.88,-12.830,-11.214,-15278.,-17828.
2064.000000000,-105.85,-12.828,-11.212,-15277.,-17828.
2065.000000000,-105.84,-12.826,-11.210,-15277.,-17827.
2066.000000000,-105.82,-12.825,-11.209,-15277.,-17827.
2067.000000000,-105.80,-12.824,-11.208,-15277.,-17827.
2068.000000000,-105.79,-12.823,-11.207,-15277.,-17827.
2069.000000000,-105.78,-12.822,-11.206,-15277.,-17827.
