time,DOLANCREEK_GAUGE,REACH_1,REACH_2,REACH_3,REACH_4,REACH_5,DEVILSRIVER
1.000000000000,-0.16051,-614.26,-2001.0,-82.210,-462.89,-8.9571,-18.641
2.000000000000,-0.16086,-637.46,-2015.0,-82.650,-463.38,-8.9618,-18.603
3.000000000000,-0.16126,-657.73,-2028.5,-83.046,-464.15,-8.9680,-18.584
4.000000000000,-0.16188,1879.9,3740.2,-53.450,-370.92,-8.9834,-18.942
5.000000000000,-0.16230,1859.6,3723.3,-53.756,-372.15,-8.9929,-18.820
6.000000000000,-0.16257,-714.14,-2073.3,-83.960,-467.04,-8.9965,-18.627
7.000000000000,-0.16281,-725.56,-2081.8,-84.184,-467.28,-9.0010,-18.601
8.000000000000,-0.16307,-736.26,-2089.3,-84.384,-467.81,-9.0058,-18.594
9.000000000000,-0.16459,1809.1,3686.1,-54.626,-375.19,-9.0555,-20.772
10.00000000000,-0.16602,1795.1,3675.5,-54.796,-377.40,-9.1026,-21.478
11.00000000000,-0.16556,-772.66,-2115.2,-84.881,-472.06,-9.0863,-19.177
12.00000000000,-0.16506,-780.38,-2118.4,-85.002,-471.73,-9.0722,-18.936
13.00000000000,-0.16479,-787.80,-2121.6,-85.109,-471.69,-9.0629,-18.832
14.00000000000,-0.16468,-795.04,-2124.4,-85.208,-471.72,-9.0577,-18.767
15.00000000000,-0.16466,-802.07,-2126.8,-85.298,-471.80,-9.0556,-18.722
16.00000000000,-0.16469,-808.62,-2128.6,-85.382,-471.94,-9.0555,-18.690
17.00000000000,-0.16470,-814.58,-2130.1,-85.459,-472.09,-9.0566,-18.667
18.00000000000,-0.16473,-819.81,-2131.4,-85.538,-472.25,-9.0585,-18.651
19.00000000000,-0.16477,-824.77,-2132.4,-85.611,-472.42,-9.0609,-18.639
20.00000000000,-0.16482,-829.53,-2133.0,-85.677,-472.58,-9.0635,-18.630
21.00000000000,-0.16488,-833.71,-2133.2,-85.735,-472.75,-9.0662,-18.624
22.00000000000,-0.16493,-837.77,-2133.2,-85.793,-472.91,-9.0690,-18.620
23.00000000000,-0.16499,-841.69,-2133.1,-85.842,-473.06,-9.0717,-18.617
24.00000000000,-0.16505,-845.39,-2133.0,-85.881,-473.21,-9.0744,-18.615
25.00000000000,-0.16510,-849.04,-2132.5,-85.919,-473.35,-9.0770,-18.614
26.00000000000,-0.16516,-852.53,-2131.8,-85.955,-473.48,-9.0795,-18.613
27.00000000000,-0.16521,-855.88,-2130.9,-85.988,-473.60,-9.0819,-18.613
28.00000000000,-0.16526,-859.21,-2129.8,-86.025,-473.70,-9.0842,-18.613
29.00000000000,-0.16532,-862.35,-2128.5,-86.060,-473.80,-9.0865,-18.613
30.00000000000,-0.16535,-865.24,-2127.2,-86.088,-473.90,-9.0886,-18.614
31.00000000000,-0.16537,-867.75,-2126.0,-86.114,-473.99,-9.0906,-18.614
32.00000000000,-0.16538,-870.10,-2124.8,-86.137,-474.07,-9.0925,-18.615
33.00000000000,-0.16538,-872.20,-2123.6,-86.158,-474.14,-9.0943,-18.615
34.00000000000,-0.16538,-873.90,-2122.4,-86.176,-474.21,-9.0960,-18.616
35.00000000000,-0.16538,-875.34,-2121.2,-86.194,-474.27,-9.0976,-18.617
36.00000000000,-0.16538,-876.73,-2119.8,-86.209,-474.33,-9.0991,-18.617
37.00000000000,-0.16538,-878.05,-2118.2,-86.223,-474.39,-9.1006,-18.618
38.00000000000,-0.16538,-879.34,-2116.7,-86.237,-474.44,-9.1019,-18.619
39.00000000000,-0.16538,-880.58,-2115.2,-86.251,-474.48,-9.1031,-18.619
40.00000000000,-0.16538,-881.77,-2113.4,-86.265,-474.52,-9.1043,-18.620
41.00000000000,-0.16538,-882.92,-2111.7,-86.277,-474.57,-9.1056,-18.635
42.00000000000,-0.16538,-884.04,-2110.0,-86.287,-474.60,-9.1066,-18.623
43.00000000000,-0.16537,-885.15,-2108.4,-86.297,-474.63,-9.1075,-18.622
44.00000000000,-0.16536,-886.16,-2106.6,-86.305,-474.65,-9.1084,-18.622
45.00000000000,-0.16536,-887.15,-2105.0,-86.310,-474.67,-9.1093,-18.623
46.00000000000,-0.16535,-888.10,-2103.5,-86.315,-474.69,-9.1101,-18.623
47.00000000000,-0.16535,-889.01,-2102.0,-86.320,-474.71,-9.1109,-18.623
48.00000000000,-0.16534,-889.80,-2100.5,-86.324,-474.72,-9.1116,-18.623
49.00000000000,-0.16534,-890.50,-2099.0,-86.329,-474.73,-9.1124,-18.623
50.00000000000,-0.16534,-891.06,-2097.6,-86.335,-474.74,-9.1131,-18.623
51.00000000000,-0.16534,-891.41,-2096.2,-86.340,-474.75,-9.1137,-18.624
52.00000000000,-0.16541,1661.9,3687.0,-56.410,-380.65,-9.1179,-18.749
53.00000000000,-0.16540,-896.56,-2098.0,-86.360,-475.22,-9.1172,-18.645
54.00000000000,-0.16537,-896.12,-2095.9,-86.362,-474.88,-9.1172,-18.636
55.00000000000,-0.16535,-895.87,-2094.1,-86.366,-474.84,-9.1173,-18.632
56.00000000000,-0.16541,1658.0,3689.4,-56.436,-380.72,-9.1210,-18.752
57.00000000000,-0.16538,-899.92,-2095.6,-86.384,-475.27,-9.1200,-18.649
58.00000000000,-0.16536,-899.01,-2093.4,-86.383,-474.92,-9.1197,-18.639
59.00000000000,-0.16534,-898.36,-2091.4,-86.385,-474.88,-9.1196,-18.635
60.00000000000,-0.16532,-897.81,-2089.7,-86.386,-474.85,-9.1197,-18.633
61.00000000000,-0.16531,-897.35,-2088.0,-86.389,-474.83,-9.1198,-18.631
62.00000000000,-0.16530,-896.94,-2086.4,-86.392,-474.82,-9.1201,-18.629
63.00000000000,-0.16529,-896.58,-2084.9,-86.395,-474.81,-9.1204,-18.628
64.00000000000,-0.16529,-896.18,-2083.4,-86.397,-474.80,-9.1207,-18.628
65.00000000000,-0.16528,-895.76,-2082.0,-86.397,-474.79,-9.1210,-18.627
66.00000000000,-0.16528,-895.40,-2080.6,-86.398,-474.79,-9.1214,-18.627
67.00000000000,-0.16527,-895.06,-2079.2,-86.398,-474.78,-9.1217,-18.626
68.00000000000,-0.16527,-894.73,-2077.8,-86.398,-474.78,-9.1221,-18.626
69.00000000000,-0.16548,1659.1,3705.4,-56.464,-380.79,-9.1310,-19.004
70.00000000000,-0.16543,-898.74,-2079.7,-86.409,-475.37,-9.1290,-18.687
71.00000000000,-0.16537,-897.80,-2077.6,-86.405,-475.00,-9.1276,-18.660
72.00000000000,-0.16534,-897.09,-2075.8,-86.404,-474.93,-9.1268,-18.649
73.00000000000,-0.16531,-896.48,-2074.2,-86.403,-474.89,-9.1264,-18.643
74.00000000000,-0.16530,-895.85,-2072.5,-86.403,-474.85,-9.1262,-18.639
75.00000000000,-0.16529,-895.28,-2070.8,-86.402,-474.82,-9.1261,-18.636
76.00000000000,-0.16528,-894.77,-2069.2,-86.401,-474.80,-9.1261,-18.633
77.00000000000,-0.16527,-894.28,-2067.7,-86.399,-474.78,-9.1263,-18.632
78.00000000000,-0.16527,-893.81,-2066.2,-86.398,-474.76,-9.1265,-18.630
79.00000000000,-0.16526,-893.35,-2064.7,-86.397,-474.75,-9.1267,-18.629
80.00000000000,-0.16526,-892.90,-2063.3,-86.395,-474.74,-9.1269,-18.628
81.00000000000,-0.16525,-892.45,-2061.9,-86.394,-474.72,-9.1272,-18.628
82.00000000000,-0.16538,1662.2,3721.2,-56.459,-380.65,-9.1328,-18.845
83.00000000000,-0.16535,-896.22,-2064.0,-86.401,-475.21,-9.1314,-18.662
84.00000000000,-0.16531,-895.08,-2062.1,-86.395,-474.85,-9.1306,-18.646
85.00000000000,-0.16529,-894.19,-2060.3,-86.392,-474.78,-9.1300,-18.640
86.00000000000,-0.16527,-893.39,-2058.7,-86.390,-474.74,-9.1296,-18.636
87.00000000000,-0.16525,-892.64,-2057.2,-86.389,-474.71,-9.1300,-18.633
88.00000000000,-0.16525,-891.93,-2055.8,-86.387,-474.68,-9.1310,-18.631
89.00000000000,-0.16524,-891.24,-2054.5,-86.386,-474.65,-9.1312,-18.630
90.00000000000,-0.16522,-890.56,-2053.1,-86.385,-474.63,-9.1313,-18.629
91.00000000000,-0.16521,-889.89,-2051.8,-86.384,-474.61,-9.1315,-18.629
92.00000000000,-0.16520,-889.23,-2050.5,-86.385,-474.59,-9.1317,-18.631
93.00000000000,-0.16574,1665.7,3732.4,-56.453,-380.85,-9.1517,-19.567
94.00000000000,-0.16561,-892.32,-2052.9,-86.398,-475.45,-9.1473,-18.792
95.00000000000,-0.16544,-890.78,-2051.0,-86.394,-475.03,-9.1430,-18.712
96.00000000000,-0.16533,-889.49,-2049.4,-86.394,-474.89,-9.1397,-18.685
97.00000000000,-0.16525,-888.34,-2047.9,-86.394,-474.78,-9.1374,-18.669
98.00000000000,-0.16520,-887.27,-2046.4,-86.395,-474.70,-9.1359,-18.657
99.00000000000,-0.16517,-886.26,-2044.9,-86.395,-474.63,-9.1349,-18.649
100.0000000000,-0.16514,-885.30,-2043.5,-86.396,-474.58,-9.1342,-18.643
101.0000000000,-0.16512,-884.36,-2042.1,-86.396,-474.53,-9.1338,-18.639
102.0000000000,-0.16510,-883.46,-2040.7,-86.397,-474.49,-9.1336,-18.635
103.0000000000,-0.16509,-882.57,-2039.4,-86.397,-474.46,-9.1334,-18.633
104.0000000000,-0.16507,-881.69,-2038.1,-86.397,-474.43,-9.1333,-18.631
105.0000000000,-0.16506,-880.82,-2036.8,-86.398,-474.40,-9.1333,-18.629
106.0000000000,-0.16505,-879.97,-2035.5,-86.398,-474.37,-9.1333,-18.628
107.0000000000,-0.16503,-879.13,-2034.3,-86.398,-474.34,-9.1332,-18.626
108.0000000000,-0.16534,1675.9,3748.6,-56.465,-380.41,-9.1451,-19.168
109.0000000000,-0.16526,-882.06,-2036.7,-86.410,-474.98,-9.1421,-18.712
110.0000000000,-0.16516,-880.49,-2034.9,-86.406,-474.58,-9.1396,-18.673
111.0000000000,-0.16510,-879.17,-2033.3,-86.406,-474.48,-9.1376,-18.658
112.0000000000,-0.16505,-877.97,-2031.8,-86.407,-474.40,-9.1362,-18.648
113.0000000000,-0.16502,-876.85,-2030.4,-86.407,-474.34,-9.1353,-18.641
114.0000000000,-0.16499,-875.78,-2029.0,-86.407,-474.29,-9.1347,-18.637
115.0000000000,-0.16497,-874.74,-2027.7,-86.407,-474.25,-9.1342,-18.633
116.0000000000,-0.16496,-873.73,-2026.5,-86.408,-474.21,-9.1339,-18.630
117.0000000000,-0.16495,-872.74,-2025.2,-86.408,-474.18,-9.1337,-18.628
118.0000000000,-0.16597,1682.4,3757.7,-56.475,-380.82,-9.1703,-20.407
119.0000000000,-0.16751,1678.7,3754.0,-56.485,-382.71,-9.2238,-21.947
120.0000000000,-0.16682,-878.59,-2030.7,-86.425,-476.93,-9.2018,-19.267
121.0000000000,-0.16613,-876.81,-2028.5,-86.422,-476.13,-9.1817,-19.002
122.0000000000,-0.16635,1678.8,3755.1,-56.489,-382.02,-9.1905,-20.034
123.0000000000,-0.16593,-878.64,-2029.7,-86.433,-476.26,-9.1745,-19.003
124.0000000000,-0.16557,-876.67,-2027.5,-86.431,-475.54,-9.1622,-18.873
125.0000000000,-0.16534,-875.06,-2025.7,-86.431,-475.17,-9.1535,-18.807
126.0000000000,-0.16519,-873.71,-2024.0,-86.430,-474.89,-9.1475,-18.762
127.0000000000,-0.16509,-872.43,-2022.3,-86.430,-474.68,-9.1435,-18.729
128.0000000000,-0.16502,-871.21,-2020.9,-86.430,-474.51,-9.1407,-18.705
129.0000000000,-0.16498,-870.04,-2019.5,-86.429,-474.38,-9.1389,-18.687
130.0000000000,-0.16528,1685.2,3763.6,-56.495,-380.39,-9.1503,-19.253
131.0000000000,-0.16560,1681.7,3760.1,-56.505,-381.07,-9.1615,-19.471
132.0000000000,-0.16540,-875.37,-2024.6,-86.444,-475.23,-9.1544,-18.822
133.0000000000,-0.16520,-873.17,-2022.3,-86.438,-474.69,-9.1485,-18.749
134.0000000000,-0.16507,-871.38,-2020.3,-86.435,-474.49,-9.1442,-18.715
135.0000000000,-0.16554,1684.4,3763.1,-56.499,-380.62,-9.1611,-19.635
136.0000000000,-0.16536,-873.00,-2021.8,-86.441,-475.11,-9.1543,-18.828
137.0000000000,-0.16517,-870.98,-2019.6,-86.435,-474.61,-9.1485,-18.749
138.0000000000,-0.16505,-869.26,-2017.7,-86.432,-474.41,-9.1442,-18.715
139.0000000000,-0.16496,-867.72,-2016.0,-86.430,-474.26,-9.1412,-18.692
140.0000000000,-0.16491,-866.31,-2014.5,-86.428,-474.15,-9.1391,-18.677
141.0000000000,-0.16487,-864.96,-2012.9,-86.426,-474.05,-9.1377,-18.665
142.0000000000,-0.16484,-863.68,-2011.5,-86.424,-473.98,-9.1367,-18.656
143.0000000000,-0.16482,-862.43,-2010.1,-86.421,-473.91,-9.1360,-18.650
144.0000000000,-0.16605,1692.9,3772.9,-56.486,-380.69,-9.1791,-20.769
145.0000000000,-0.16586,1689.5,3769.3,-56.494,-381.25,-9.1735,-19.156
146.0000000000,-0.16742,1686.6,3766.3,-56.499,-382.66,-9.2296,-22.168
147.0000000000,-0.16673,-870.14,-2018.0,-86.437,-476.80,-9.2060,-19.312
148.0000000000,-0.16603,-867.99,-2015.5,-86.434,-475.95,-9.1849,-19.034
149.0000000000,-0.16585,1688.1,3768.2,-56.502,-381.48,-9.1795,-19.381
150.0000000000,-0.16551,-869.16,-2016.5,-86.447,-475.65,-9.1659,-18.920
151.0000000000,-0.16525,-866.97,-2014.3,-86.445,-474.97,-9.1565,-18.832
152.0000000000,-0.16509,-865.15,-2012.3,-86.445,-474.66,-9.1499,-18.781
153.0000000000,-0.16498,-863.56,-2010.5,-86.444,-474.42,-9.1454,-18.745
154.0000000000,-0.16495,1692.1,3772.8,-56.511,-380.12,-9.1448,-18.789
155.0000000000,-0.16490,-865.32,-2012.1,-86.455,-474.54,-9.1417,-18.711
156.0000000000,-0.16485,-863.27,-2010.0,-86.450,-474.09,-9.1398,-18.691
157.0000000000,-0.16482,-861.51,-2008.1,-86.448,-473.97,-9.1385,-18.677
158.0000000000,-0.16480,-859.91,-2006.4,-86.446,-473.89,-9.1379,-18.685
159.0000000000,-0.16522,1695.7,3776.8,-56.511,-380.01,-9.1532,-19.413
160.0000000000,-0.16511,-861.72,-2008.3,-86.454,-474.55,-9.1487,-18.776
161.0000000000,-0.16497,-859.72,-2006.2,-86.450,-474.11,-9.1448,-18.719
162.0000000000,-0.16488,-857.99,-2004.4,-86.448,-473.97,-9.1417,-18.693
163.0000000000,-0.16482,-856.52,-2002.8,-86.447,-473.86,-9.1395,-18.677
164.0000000000,-0.16478,-855.13,-2001.3,-86.446,-473.77,-9.1381,-18.666
165.0000000000,-0.16503,1700.4,3781.8,-56.510,-379.77,-9.1476,-19.136
166.0000000000,-0.16743,1697.1,3778.4,-56.519,-382.12,-9.2304,-22.982
167.0000000000,-0.16698,1694.2,3775.4,-56.524,-382.50,-9.2162,-19.688
168.0000000000,-0.16619,-862.59,-2008.8,-86.464,-476.29,-9.1928,-19.101
169.0000000000,-0.16584,1694.1,3775.5,-56.527,-381.40,-9.1822,-19.271
170.0000000000,-0.16552,1691.5,3772.7,-56.540,-381.39,-9.1705,-19.013
171.0000000000,-0.16525,-864.82,-2011.3,-86.479,-475.25,-9.1593,-18.854
172.0000000000,-0.16506,-862.04,-2008.4,-86.474,-474.59,-9.1519,-18.796
173.0000000000,-0.16494,-859.79,-2006.1,-86.473,-474.31,-9.1469,-18.757
174.0000000000,-0.16487,-857.79,-2004.1,-86.472,-474.11,-9.1435,-18.729
175.0000000000,-0.16481,-855.97,-2002.2,-86.471,-473.95,-9.1411,-18.708
176.0000000000,-0.16478,-854.28,-2000.4,-86.470,-473.83,-9.1395,-18.692
177.0000000000,-0.16475,-852.67,-1998.7,-86.468,-473.73,-9.1383,-18.679
178.0000000000,-0.16473,-851.17,-1997.1,-86.467,-473.65,-9.1375,-18.670
179.0000000000,-0.16471,-849.74,-1995.6,-86.465,-473.59,-9.1368,-18.662
180.0000000000,-0.16470,-848.35,-1994.2,-86.464,-473.54,-9.1364,-18.657
181.0000000000,-0.16531,1707.1,3788.9,-56.529,-379.82,-9.1582,-19.709
182.0000000000,-0.16517,-850.39,-1996.3,-86.472,-474.41,-9.1529,-18.830
183.0000000000,-0.16513,1705.7,3787.3,-56.534,-379.91,-9.1536,-18.979
184.0000000000,-0.16498,-851.45,-1997.5,-86.476,-474.32,-9.1478,-18.749
185.0000000000,-0.16486,-849.22,-1995.4,-86.470,-473.85,-9.1439,-18.712
186.0000000000,-0.16479,-847.35,-1993.5,-86.468,-473.70,-9.1410,-18.692
187.0000000000,-0.16474,-845.70,-1991.8,-86.466,-473.59,-9.1391,-18.678
188.0000000000,-0.16471,-844.17,-1990.2,-86.464,-473.50,-9.1377,-18.668
189.0000000000,-0.16468,-842.73,-1988.7,-86.462,-473.44,-9.1367,-18.660
190.0000000000,-0.16467,-841.38,-1987.3,-86.461,-473.38,-9.1360,-18.655
191.0000000000,-0.16465,-840.07,-1985.9,-86.459,-473.34,-9.1355,-18.650
192.0000000000,-0.16464,-838.80,-1984.6,-86.458,-473.30,-9.1351,-18.647
193.0000000000,-0.16463,-837.57,-1983.3,-86.456,-473.26,-9.1348,-18.644
194.0000000000,-0.16463,-836.37,-1982.1,-86.454,-473.23,-9.1345,-18.642
195.0000000000,-0.16462,-835.18,-1980.9,-86.453,-473.20,-9.1343,-18.640
196.0000000000,-0.16477,1720.1,3802.0,-56.519,-379.14,-9.1406,-18.907
197.0000000000,-0.16635,1716.6,3798.3,-56.528,-380.83,-9.1952,-21.455
198.0000000000,-0.16681,1713.8,3795.2,-56.534,-381.69,-9.2115,-20.569
199.0000000000,-0.16630,1711.2,3792.6,-56.540,-381.67,-9.1973,-19.406
200.0000000000,-0.16598,1708.9,3790.1,-56.546,-381.50,-9.1881,-19.437
201.0000000000,-0.16553,-847.40,-1993.7,-86.486,-475.29,-9.1717,-18.963
202.0000000000,-0.16526,1709.6,3790.9,-56.549,-380.41,-9.1625,-18.935
203.0000000000,-0.16512,1707.2,3788.4,-56.559,-380.51,-9.1568,-18.933
204.0000000000,-0.16497,-848.95,-1995.5,-86.499,-474.47,-9.1495,-18.788
205.0000000000,-0.16486,-846.06,-1992.5,-86.495,-473.90,-9.1449,-18.748
206.0000000000,-0.16479,-843.70,-1990.0,-86.494,-473.68,-9.1416,-18.721
207.0000000000,-0.16474,-841.64,-1987.8,-86.493,-473.53,-9.1394,-18.702
208.0000000000,-0.16478,1714.4,3795.8,-56.559,-379.31,-9.1413,-18.811
209.0000000000,-0.16475,-842.69,-1988.9,-86.502,-473.78,-9.1389,-18.696
210.0000000000,-0.16495,1713.8,3795.1,-56.564,-379.40,-9.1467,-19.091
211.0000000000,-0.16488,-843.03,-1989.4,-86.506,-473.88,-9.1431,-18.735
212.0000000000,-0.16479,-840.54,-1986.8,-86.501,-473.44,-9.1404,-18.698
213.0000000000,-0.16474,-838.45,-1984.6,-86.499,-473.32,-9.1383,-18.681
214.0000000000,-0.16471,-836.57,-1982.7,-86.497,-473.23,-9.1370,-18.676
215.0000000000,-0.16468,-834.84,-1980.8,-86.494,-473.15,-9.1359,-18.663
216.0000000000,-0.16466,-833.22,-1979.1,-86.492,-473.09,-9.1351,-18.656
217.0000000000,-0.16465,-831.67,-1977.5,-86.490,-473.04,-9.1345,-18.651
218.0000000000,-0.16464,-830.19,-1976.0,-86.487,-473.00,-9.1341,-18.648
219.0000000000,-0.16464,-828.79,-1974.5,-86.485,-472.96,-9.1338,-18.645
220.0000000000,-0.16463,-827.41,-1973.1,-86.481,-472.93,-9.1335,-18.642
221.0000000000,-0.16463,-826.13,-1971.7,-86.478,-472.90,-9.1333,-18.641
222.0000000000,-0.16462,-824.85,-1970.4,-86.475,-472.87,-9.1331,-18.639
223.0000000000,-0.16463,-823.60,-1969.1,-86.471,-472.86,-9.1334,-18.662
224.0000000000,-0.16470,1731.8,3813.8,-56.534,-378.73,-9.1368,-18.775
225.0000000000,-0.16468,-825.87,-1971.5,-86.474,-473.28,-9.1353,-18.660
226.0000000000,-0.16465,-824.01,-1969.7,-86.467,-472.91,-9.1344,-18.649
227.0000000000,-0.16464,-822.42,-1968.1,-86.463,-472.85,-9.1336,-18.644
228.0000000000,-0.16462,-820.97,-1966.6,-86.459,-472.80,-9.1331,-18.642
229.0000000000,-0.16461,-819.61,-1965.2,-86.456,-472.77,-9.1327,-18.639
230.0000000000,-0.16461,-818.31,-1963.9,-86.452,-472.73,-9.1324,-18.637
231.0000000000,-0.16460,-817.06,-1962.6,-86.448,-472.71,-9.1322,-18.637
232.0000000000,-0.16460,-815.85,-1961.4,-86.445,-472.68,-9.1319,-18.634
233.0000000000,-0.16459,-814.66,-1960.1,-86.441,-472.65,-9.1317,-18.633
234.0000000000,-0.16464,1740.7,3822.7,-56.504,-378.50,-9.1342,-18.717
235.0000000000,-0.16462,-817.01,-1962.7,-86.444,-473.05,-9.1330,-18.646
236.0000000000,-0.16590,1739.0,3820.7,-56.503,-379.57,-9.1779,-20.859
237.0000000000,-0.16563,1735.8,3817.3,-56.508,-380.05,-9.1692,-19.042
238.0000000000,-0.16545,1733.3,3814.5,-56.510,-380.05,-9.1653,-19.161
239.0000000000,-0.16683,1731.0,3811.9,-56.512,-381.20,-9.2132,-21.693
240.0000000000,-0.16761,1729.0,3809.6,-56.514,-382.25,-9.2405,-21.552
241.0000000000,-0.16672,-827.43,-1974.2,-86.452,-476.13,-9.2115,-19.354
242.0000000000,-0.16596,-824.83,-1971.2,-86.448,-475.14,-9.1872,-19.087
243.0000000000,-0.16547,-822.54,-1968.8,-86.448,-474.52,-9.1696,-18.960
244.0000000000,-0.16517,-820.61,-1966.7,-86.446,-474.05,-9.1575,-18.876
245.0000000000,-0.16499,-818.88,-1964.9,-86.444,-473.70,-9.1494,-18.818
246.0000000000,-0.16545,1736.9,3818.4,-56.509,-379.73,-9.1652,-19.782
247.0000000000,-0.16524,-820.37,-1966.4,-86.451,-474.14,-9.1564,-18.904
248.0000000000,-0.16549,1736.0,3817.4,-56.511,-379.77,-9.1660,-19.595
249.0000000000,-0.16553,1733.2,3814.5,-56.518,-380.18,-9.1672,-19.368
250.0000000000,-0.16525,-823.29,-1969.7,-86.455,-474.18,-9.1570,-18.878
251.0000000000,-0.16503,-820.62,-1967.0,-86.448,-473.56,-9.1494,-18.801
252.0000000000,-0.16526,1735.7,3816.9,-56.511,-379.43,-9.1577,-19.397
253.0000000000,-0.16516,1732.9,3814.1,-56.518,-379.71,-9.1535,-18.939
254.0000000000,-0.16517,1730.7,3811.6,-56.522,-379.73,-9.1541,-19.100
255.0000000000,-0.16501,-825.36,-1972.1,-86.459,-473.76,-9.1474,-18.796
256.0000000000,-0.16488,-822.41,-1969.2,-86.453,-473.21,-9.1426,-18.744
257.0000000000,-0.16479,-820.00,-1966.7,-86.449,-473.02,-9.1392,-18.717
258.0000000000,-0.16474,-817.95,-1964.5,-86.446,-472.87,-9.1367,-18.698
259.0000000000,-0.16470,-816.13,-1962.5,-86.443,-472.76,-9.1350,-18.684
260.0000000000,-0.16499,1739.7,3820.9,-56.507,-378.76,-9.1456,-19.216
261.0000000000,-0.16552,1736.6,3817.7,-56.514,-379.61,-9.1639,-19.812
262.0000000000,-0.16543,1734.1,3815.1,-56.518,-379.75,-9.1615,-19.126
263.0000000000,-0.16885,1732.0,3812.8,-56.520,-382.57,-9.2803,-25.155
264.0000000000,-0.17084,1729.1,3810.5,-56.527,-385.16,-9.3500,-24.923
265.0000000000,-0.16903,-828.08,-1973.5,-86.480,-478.96,-9.2938,-20.110
266.0000000000,-0.16746,-826.03,-1971.1,-86.491,-477.47,-9.2452,-19.551
267.0000000000,-0.16646,-824.04,-1968.7,-86.498,-476.34,-9.2097,-19.293
268.0000000000,-0.16584,-822.08,-1966.4,-86.500,-475.46,-9.1853,-19.126
269.0000000000,-0.16546,-820.22,-1964.4,-86.498,-474.79,-9.1690,-19.008
270.0000000000,-0.16521,-818.54,-1962.5,-86.501,-474.29,-9.1582,-18.923
271.0000000000,-0.16506,-817.36,-1960.7,-86.501,-473.90,-9.1509,-18.860
272.0000000000,-0.16546,1738.2,3822.7,-56.567,-379.84,-9.1642,-19.675
273.0000000000,-0.16528,-819.41,-1962.3,-86.510,-474.22,-9.1563,-18.916
274.0000000000,-0.16509,-817.47,-1960.1,-86.505,-473.65,-9.1499,-18.826
275.0000000000,-0.16497,-815.84,-1958.3,-86.505,-473.40,-9.1453,-18.782
276.0000000000,-0.16489,-814.43,-1956.6,-86.504,-473.22,-9.1419,-18.752
277.0000000000,-0.16483,-813.15,-1955.0,-86.503,-473.07,-9.1395,-18.729
278.0000000000,-0.16479,-811.86,-1953.6,-86.502,-472.95,-9.1378,-18.713
279.0000000000,-0.16477,-810.55,-1952.2,-86.502,-472.86,-9.1368,-18.708
280.0000000000,-0.16475,-809.34,-1950.9,-86.503,-472.79,-9.1358,-18.691
281.0000000000,-0.16474,-808.13,-1949.6,-86.505,-472.72,-9.1351,-18.683
282.0000000000,-0.16473,-807.02,-1948.4,-86.508,-472.67,-9.1345,-18.676
283.0000000000,-0.16474,-805.91,-1947.1,-86.511,-472.62,-9.1341,-18.672
284.0000000000,-0.16474,-804.83,-1945.9,-86.515,-472.58,-9.1337,-18.668
285.0000000000,-0.16474,-803.79,-1944.6,-86.516,-472.55,-9.1334,-18.664
286.0000000000,-0.16476,-802.75,-1943.4,-86.518,-472.53,-9.1336,-18.685
287.0000000000,-0.16522,1752.6,3839.4,-56.586,-378.71,-9.1500,-19.436
288.0000000000,-0.16594,1749.0,3835.6,-56.598,-379.78,-9.1750,-20.189
289.0000000000,-0.16813,1746.1,3832.5,-56.605,-381.83,-9.2512,-23.222
290.0000000000,-0.16733,1743.3,3829.5,-56.610,-381.96,-9.2261,-19.618
291.0000000000,-0.16643,-813.59,-1954.7,-86.549,-475.59,-9.1985,-19.173
292.0000000000,-0.16585,-811.03,-1952.2,-86.547,-474.64,-9.1784,-19.038
293.0000000000,-0.16548,-808.92,-1950.1,-86.545,-474.11,-9.1642,-18.925
294.0000000000,-0.16525,-807.12,-1948.4,-86.544,-473.72,-9.1546,-18.858
295.0000000000,-0.16511,-805.54,-1946.8,-86.543,-473.43,-9.1482,-18.809
296.0000000000,-0.16501,-804.03,-1945.4,-86.543,-473.20,-9.1438,-18.774
297.0000000000,-0.16495,-802.59,-1943.9,-86.541,-473.03,-9.1408,-18.747
298.0000000000,-0.16491,-801.21,-1942.5,-86.538,-472.89,-9.1387,-18.727
299.0000000000,-0.16488,-799.94,-1941.1,-86.536,-472.78,-9.1372,-18.711
300.0000000000,-0.16486,-798.71,-1939.8,-86.533,-472.69,-9.1360,-18.699
301.0000000000,-0.16484,-797.52,-1938.5,-86.530,-472.62,-9.1352,-18.690
302.0000000000,-0.16483,-796.33,-1937.3,-86.528,-472.56,-9.1346,-18.683
303.0000000000,-0.16482,-795.09,-1936.2,-86.525,-472.51,-9.1340,-18.677
304.0000000000,-0.16483,1760.5,3846.6,-56.589,-378.32,-9.1353,-18.709
305.0000000000,-0.16483,-797.20,-1938.8,-86.530,-472.84,-9.1341,-18.675
306.0000000000,-0.16481,-795.27,-1937.0,-86.524,-472.48,-9.1335,-18.670
307.0000000000,-0.16481,-793.63,-1935.5,-86.521,-472.41,-9.1331,-18.666
308.0000000000,-0.16512,1762.1,3847.4,-56.587,-378.47,-9.1448,-19.217
309.0000000000,-0.16514,1758.8,3843.7,-56.596,-378.94,-9.1455,-18.906
310.0000000000,-0.16530,1756.0,3840.6,-56.601,-379.16,-9.1516,-19.200
311.0000000000,-0.16538,1753.7,3837.9,-56.605,-379.31,-9.1546,-19.166
312.0000000000,-0.16520,-802.63,-1946.2,-86.542,-473.40,-9.1478,-18.797
313.0000000000,-0.16531,1754.5,3838.2,-56.601,-378.93,-9.1527,-19.193
314.0000000000,-0.16516,-802.16,-1946.1,-86.542,-473.33,-9.1463,-18.793
315.0000000000,-0.16503,-799.46,-1943.5,-86.536,-472.85,-9.1418,-18.744
316.0000000000,-0.16499,1757.1,3840.3,-56.598,-378.55,-9.1412,-18.812
317.0000000000,-0.16494,-799.88,-1944.3,-86.539,-473.01,-9.1381,-18.741
318.0000000000,-0.16489,-797.41,-1942.0,-86.531,-472.58,-9.1358,-18.704
319.0000000000,-0.16485,-795.32,-1939.9,-86.526,-472.46,-9.1341,-18.690
320.0000000000,-0.16482,-793.43,-1938.1,-86.522,-472.38,-9.1329,-18.681
321.0000000000,-0.16480,-791.66,-1936.4,-86.517,-472.31,-9.1319,-18.674
322.0000000000,-0.16479,-789.96,-1934.9,-86.513,-472.26,-9.1312,-18.669
323.0000000000,-0.16478,-788.34,-1933.4,-86.508,-472.21,-9.1306,-18.665
324.0000000000,-0.16477,-786.80,-1932.0,-86.503,-472.17,-9.1302,-18.662
325.0000000000,-0.16476,-785.34,-1930.6,-86.499,-472.14,-9.1298,-18.659
326.0000000000,-0.16486,1770.4,3852.3,-56.561,-378.03,-9.1340,-18.833
327.0000000000,-0.16493,1767.1,3848.6,-56.566,-378.48,-9.1365,-18.854
328.0000000000,-0.16554,1764.5,3845.5,-56.568,-379.05,-9.1578,-19.837
329.0000000000,-0.16588,1762.2,3842.8,-56.570,-379.53,-9.1698,-19.776
330.0000000000,-0.16556,-793.99,-1941.3,-86.505,-473.64,-9.1590,-18.939
331.0000000000,-0.16527,-791.03,-1938.6,-86.496,-473.04,-9.1497,-18.820
332.0000000000,-0.16508,-788.62,-1936.4,-86.491,-472.77,-9.1428,-18.771
333.0000000000,-0.16496,-786.55,-1934.5,-86.486,-472.58,-9.1381,-18.740
334.0000000000,-0.16489,-784.66,-1932.8,-86.481,-472.42,-9.1348,-18.718
335.0000000000,-0.16483,-782.89,-1931.2,-86.477,-472.31,-9.1325,-18.701
336.0000000000,-0.16480,-781.25,-1929.7,-86.472,-472.21,-9.1309,-18.689
337.0000000000,-0.16477,-779.68,-1928.3,-86.466,-472.14,-9.1296,-18.680
338.0000000000,-0.16475,-778.17,-1926.9,-86.461,-472.07,-9.1287,-18.672
339.0000000000,-0.16473,-776.71,-1925.6,-86.454,-472.02,-9.1280,-18.667
340.0000000000,-0.16485,1779.0,3857.3,-56.514,-377.92,-9.1328,-18.881
341.0000000000,-0.16481,-778.60,-1928.1,-86.453,-472.45,-9.1307,-18.696
342.0000000000,-0.16476,-776.57,-1926.3,-86.443,-472.08,-9.1293,-18.676
343.0000000000,-0.16474,-774.83,-1924.8,-86.437,-472.00,-9.1281,-18.668
344.0000000000,-0.16471,-773.24,-1923.4,-86.431,-471.94,-9.1273,-18.663
345.0000000000,-0.16470,-771.76,-1922.1,-86.426,-471.90,-9.1266,-18.658
346.0000000000,-0.16469,-770.37,-1920.8,-86.421,-471.86,-9.1260,-18.655
347.0000000000,-0.16467,-769.05,-1919.6,-86.415,-471.83,-9.1255,-18.653
348.0000000000,-0.16466,-767.76,-1918.5,-86.409,-471.80,-9.1251,-18.651
349.0000000000,-0.16465,-766.50,-1917.4,-86.403,-471.77,-9.1247,-18.649
350.0000000000,-0.16464,-765.26,-1916.3,-86.396,-471.75,-9.1244,-18.648
351.0000000000,-0.16463,-764.05,-1915.2,-86.389,-471.73,-9.1240,-18.647
352.0000000000,-0.16462,-762.86,-1914.2,-86.383,-471.70,-9.1237,-18.646
353.0000000000,-0.16461,-761.71,-1913.2,-86.377,-471.68,-9.1234,-18.645
354.0000000000,-0.16460,-760.58,-1912.2,-86.371,-471.66,-9.1231,-18.644
355.0000000000,-0.16508,1794.9,3870.5,-56.431,-377.88,-9.1408,-19.484
356.0000000000,-0.16515,1791.3,3866.5,-56.435,-378.45,-9.1436,-19.095
357.0000000000,-0.16497,-765.94,-1918.4,-86.370,-472.61,-9.1373,-18.768
358.0000000000,-0.16482,-763.77,-1916.3,-86.359,-472.14,-9.1327,-18.723
359.0000000000,-0.16472,-761.98,-1914.6,-86.353,-471.99,-9.1292,-18.700
360.0000000000,-0.16482,1793.9,3868.5,-56.413,-377.83,-9.1332,-18.964
361.0000000000,-0.16508,1790.7,3865.0,-56.417,-378.42,-9.1419,-19.283
362.0000000000,-0.16521,1788.1,3862.0,-56.418,-378.65,-9.1468,-19.272
363.0000000000,-0.16501,-768.52,-1922.2,-86.352,-472.76,-9.1394,-18.806
364.0000000000,-0.16484,-765.88,-1919.7,-86.341,-472.23,-9.1337,-18.746
365.0000000000,-0.16473,-763.74,-1917.6,-86.334,-472.04,-9.1296,-18.717
366.0000000000,-0.16466,-761.91,-1915.7,-86.328,-471.90,-9.1266,-18.697
367.0000000000,-0.16461,-760.29,-1914.0,-86.322,-471.79,-9.1245,-18.683
368.0000000000,-0.16458,-758.78,-1912.5,-86.316,-471.71,-9.1230,-18.673
369.0000000000,-0.16456,-757.35,-1911.0,-86.310,-471.64,-9.1219,-18.665
370.0000000000,-0.16454,-756.00,-1909.6,-86.305,-471.59,-9.1210,-18.659
371.0000000000,-0.16453,-754.70,-1908.3,-86.298,-471.54,-9.1203,-18.654
372.0000000000,-0.16452,-753.44,-1907.1,-86.292,-471.50,-9.1198,-18.650
373.0000000000,-0.16451,-752.24,-1905.9,-86.286,-471.47,-9.1193,-18.647
374.0000000000,-0.16451,-751.06,-1904.7,-86.280,-471.44,-9.1189,-18.645
375.0000000000,-0.16450,-749.92,-1903.6,-86.274,-471.41,-9.1185,-18.643
376.0000000000,-0.16449,-748.78,-1902.5,-86.268,-471.38,-9.1181,-18.641
377.0000000000,-0.16449,-747.66,-1901.5,-86.261,-471.36,-9.1178,-18.640
378.0000000000,-0.16448,-746.54,-1900.4,-86.255,-471.33,-9.1175,-18.638
379.0000000000,-0.16448,-745.46,-1899.4,-86.249,-471.31,-9.1172,-18.637
380.0000000000,-0.16447,-744.40,-1898.4,-86.243,-471.29,-9.1169,-18.636
381.0000000000,-0.16447,-743.36,-1897.4,-86.236,-471.28,-9.1166,-18.636
382.0000000000,-0.16446,-742.34,-1896.4,-86.230,-471.26,-9.1163,-18.635
383.0000000000,-0.16446,-741.34,-1895.4,-86.223,-471.24,-9.1160,-18.634
384.0000000000,-0.16445,-740.35,-1894.5,-86.217,-471.22,-9.1158,-18.634
385.0000000000,-0.16445,-739.37,-1893.6,-86.211,-471.21,-9.1155,-18.633
386.0000000000,-0.16444,-738.40,-1892.6,-86.204,-471.19,-9.1152,-18.632
387.0000000000,-0.16444,-737.45,-1891.7,-86.198,-471.17,-9.1150,-18.632
388.0000000000,-0.16443,-736.51,-1890.9,-86.192,-471.16,-9.1147,-18.631
389.0000000000,-0.16447,1818.8,3891.6,-56.253,-377.01,-9.1170,-18.704
390.0000000000,-0.16446,-739.34,-1894.0,-86.191,-471.56,-9.1157,-18.643
391.0000000000,-0.16444,-737.74,-1892.5,-86.182,-471.21,-9.1150,-18.637
392.0000000000,-0.16443,-736.41,-1891.2,-86.175,-471.16,-9.1145,-18.635
393.0000000000,-0.16442,-735.21,-1890.0,-86.169,-471.13,-9.1140,-18.633
394.0000000000,-0.16441,-734.16,-1888.9,-86.162,-471.10,-9.1136,-18.631
395.0000000000,-0.16441,-733.19,-1887.9,-86.156,-471.07,-9.1132,-18.630
396.0000000000,-0.16440,-732.25,-1886.9,-86.150,-471.05,-9.1129,-18.629
397.0000000000,-0.16440,-731.35,-1885.9,-86.144,-471.03,-9.1126,-18.628
398.0000000000,-0.16439,-730.45,-1884.9,-86.137,-471.01,-9.1123,-18.628
399.0000000000,-0.16439,-729.57,-1883.9,-86.131,-470.99,-9.1120,-18.630
400.0000000000,-0.16438,-728.69,-1883.0,-86.125,-470.98,-9.1117,-18.627
401.0000000000,-0.16437,-727.85,-1882.0,-86.119,-470.96,-9.1114,-18.626
402.0000000000,-0.16437,-727.02,-1881.1,-86.112,-470.94,-9.1112,-18.625
403.0000000000,-0.16437,-726.20,-1880.2,-86.106,-470.93,-9.1109,-18.625
404.0000000000,-0.16436,-725.40,-1879.3,-86.100,-470.91,-9.1106,-18.624
405.0000000000,-0.16436,-724.60,-1878.4,-86.094,-470.89,-9.1104,-18.624
406.0000000000,-0.16435,-723.81,-1877.6,-86.088,-470.88,-9.1101,-18.623
407.0000000000,-0.16435,-723.02,-1876.7,-86.083,-470.86,-9.1099,-18.623
408.0000000000,-0.16435,-722.25,-1875.8,-86.077,-470.85,-9.1096,-18.622
409.0000000000,-0.16434,-721.48,-1875.0,-86.070,-470.83,-9.1093,-18.622
410.0000000000,-0.16434,-720.72,-1874.1,-86.064,-470.81,-9.1091,-18.621
411.0000000000,-0.16433,-719.97,-1873.3,-86.058,-470.80,-9.1088,-18.621
412.0000000000,-0.16433,-719.23,-1872.5,-86.052,-470.78,-9.1086,-18.621
413.0000000000,-0.16433,-718.50,-1871.6,-86.046,-470.77,-9.1083,-18.620
414.0000000000,-0.16432,-717.77,-1870.8,-86.039,-470.75,-9.1081,-18.620
415.0000000000,-0.16432,-717.05,-1870.0,-86.033,-470.74,-9.1078,-18.619
416.0000000000,-0.16431,-716.34,-1869.2,-86.026,-470.72,-9.1076,-18.619
417.0000000000,-0.16431,-715.62,-1868.4,-86.020,-470.71,-9.1074,-18.618
418.0000000000,-0.16430,-714.91,-1867.6,-86.013,-470.69,-9.1071,-18.618
419.0000000000,-0.16430,-714.21,-1866.8,-86.007,-470.68,-9.1069,-18.617
420.0000000000,-0.16429,-713.51,-1866.0,-86.001,-470.66,-9.1066,-18.617
421.0000000000,-0.16432,1842.2,3916.4,-56.061,-376.50,-9.1084,-18.667
422.0000000000,-0.16473,1838.5,3912.2,-56.066,-377.23,-9.1229,-19.356
423.0000000000,-0.16476,1835.4,3908.7,-56.066,-377.43,-9.1241,-18.963
424.0000000000,-0.16460,-722.22,-1876.0,-86.000,-471.56,-9.1185,-18.721
425.0000000000,-0.16449,-720.21,-1873.8,-85.990,-471.09,-9.1146,-18.684
426.0000000000,-0.16442,-718.64,-1872.1,-85.983,-470.96,-9.1120,-18.685
427.0000000000,-0.16436,-717.30,-1870.6,-85.977,-470.86,-9.1098,-18.655
428.0000000000,-0.16433,-716.11,-1869.2,-85.971,-470.78,-9.1082,-18.646
429.0000000000,-0.16430,-715.02,-1867.9,-85.965,-470.72,-9.1070,-18.637
430.0000000000,-0.16428,-714.00,-1866.7,-85.959,-470.66,-9.1061,-18.631
431.0000000000,-0.16427,-713.04,-1865.6,-85.953,-470.62,-9.1054,-18.627
432.0000000000,-0.16426,-712.13,-1864.5,-85.947,-470.59,-9.1048,-18.623
433.0000000000,-0.16425,-711.24,-1863.5,-85.941,-470.56,-9.1044,-18.621
434.0000000000,-0.16426,1844.6,3919.1,-56.001,-376.38,-9.1056,-18.650
435.0000000000,-0.16425,-713.91,-1866.4,-85.939,-470.92,-9.1044,-18.623
436.0000000000,-0.16424,-712.44,-1864.8,-85.929,-470.57,-9.1039,-18.619
437.0000000000,-0.16423,-711.24,-1863.5,-85.923,-470.51,-9.1034,-18.617
438.0000000000,-0.16422,-710.18,-1862.2,-85.917,-470.48,-9.1030,-18.615
439.0000000000,-0.16421,-709.20,-1861.1,-85.911,-470.45,-9.1026,-18.614
440.0000000000,-0.16421,-708.27,-1860.0,-85.905,-470.43,-9.1023,-18.613
441.0000000000,-0.16420,-707.39,-1859.0,-85.899,-470.41,-9.1020,-18.612
442.0000000000,-0.16419,-706.55,-1858.0,-85.893,-470.39,-9.1017,-18.611
443.0000000000,-0.16419,-705.73,-1857.0,-85.887,-470.37,-9.1014,-18.610
444.0000000000,-0.16418,-704.93,-1856.0,-85.880,-470.35,-9.1012,-18.609
445.0000000000,-0.16418,-704.17,-1855.1,-85.874,-470.33,-9.1009,-18.609
446.0000000000,-0.16417,-703.41,-1854.2,-85.868,-470.32,-9.1007,-18.608
447.0000000000,-0.16417,-702.67,-1853.2,-85.862,-470.30,-9.1004,-18.608
448.0000000000,-0.16426,1853.1,3929.3,-55.923,-376.19,-9.1044,-18.772
449.0000000000,-0.16423,-705.59,-1856.4,-85.861,-470.75,-9.1028,-18.634
450.0000000000,-0.16420,-704.23,-1854.9,-85.851,-470.39,-9.1018,-18.622
451.0000000000,-0.16420,1851.9,3928.0,-55.912,-376.18,-9.1025,-18.645
452.0000000000,-0.16418,-706.50,-1857.3,-85.850,-470.71,-9.1010,-18.619
453.0000000000,-0.16416,-704.94,-1855.6,-85.840,-470.35,-9.1003,-18.614
454.0000000000,-0.16415,-703.68,-1854.1,-85.834,-470.29,-9.0997,-18.611
455.0000000000,-0.16414,-702.58,-1852.8,-85.828,-470.25,-9.0992,-18.609
456.0000000000,-0.16413,-701.56,-1851.6,-85.823,-470.22,-9.0988,-18.608
457.0000000000,-0.16412,-700.61,-1850.5,-85.817,-470.20,-9.0984,-18.606
458.0000000000,-0.16411,-699.71,-1849.4,-85.811,-470.17,-9.0981,-18.605
459.0000000000,-0.16447,1856.2,3933.3,-55.872,-376.28,-9.1112,-19.221
460.0000000000,-0.16438,-702.37,-1852.3,-85.810,-470.85,-9.1075,-18.703
461.0000000000,-0.16430,1854.1,3931.0,-55.867,-376.31,-9.1061,-18.687
462.0000000000,-0.16423,-704.08,-1854.2,-85.805,-470.77,-9.1029,-18.651
463.0000000000,-0.16422,1852.6,3929.3,-55.862,-376.23,-9.1032,-18.703
464.0000000000,-0.16418,-705.36,-1855.7,-85.800,-470.71,-9.1008,-18.637
465.0000000000,-0.16414,-703.50,-1853.6,-85.790,-470.31,-9.0993,-18.626
466.0000000000,-0.16412,-701.99,-1851.9,-85.784,-470.22,-9.0982,-18.619
467.0000000000,-0.16409,-700.68,-1850.4,-85.778,-470.16,-9.0973,-18.614
468.0000000000,-0.16407,-699.49,-1849.2,-85.773,-470.12,-9.0967,-18.611
469.0000000000,-0.16406,-698.39,-1848.1,-85.767,-470.09,-9.0963,-18.617
470.0000000000,-0.16405,-697.36,-1847.0,-85.761,-470.05,-9.0958,-18.607
471.0000000000,-0.16404,-696.39,-1846.0,-85.755,-470.03,-9.0954,-18.604
472.0000000000,-0.16403,-695.45,-1845.0,-85.750,-470.00,-9.0950,-18.603
473.0000000000,-0.16401,-694.56,-1844.1,-85.744,-469.98,-9.0947,-18.601
474.0000000000,-0.16400,-693.69,-1843.2,-85.738,-469.96,-9.0944,-18.600
475.0000000000,-0.16404,1862.2,3940.2,-55.799,-375.81,-9.0967,-18.678
476.0000000000,-0.16402,-696.43,-1846.1,-85.737,-470.36,-9.0954,-18.612
477.0000000000,-0.16400,-694.96,-1844.7,-85.727,-470.01,-9.0947,-18.605
478.0000000000,-0.16398,-693.77,-1843.4,-85.721,-469.95,-9.0941,-18.602
479.0000000000,-0.16397,-692.71,-1842.4,-85.715,-469.92,-9.0936,-18.600
480.0000000000,-0.16396,-691.74,-1841.4,-85.709,-469.89,-9.0932,-18.599
481.0000000000,-0.16395,-690.83,-1840.4,-85.702,-469.86,-9.0928,-18.598
482.0000000000,-0.16394,-689.96,-1839.5,-85.696,-469.84,-9.0925,-18.597
483.0000000000,-0.16393,-689.13,-1838.6,-85.690,-469.82,-9.0922,-18.596
484.0000000000,-0.16392,-688.31,-1837.8,-85.684,-469.80,-9.0919,-18.595
485.0000000000,-0.16391,-687.52,-1837.0,-85.678,-469.78,-9.0917,-18.594
486.0000000000,-0.16390,-686.74,-1836.2,-85.672,-469.77,-9.0914,-18.594
487.0000000000,-0.16389,-685.99,-1835.4,-85.666,-469.75,-9.0912,-18.593
488.0000000000,-0.16388,-685.26,-1834.6,-85.660,-469.73,-9.0909,-18.593
489.0000000000,-0.16387,-684.53,-1833.9,-85.654,-469.72,-9.0907,-18.592
490.0000000000,-0.16387,-683.82,-1833.1,-85.648,-469.70,-9.0905,-18.592
491.0000000000,-0.16386,-683.12,-1832.4,-85.642,-469.69,-9.0902,-18.591
492.0000000000,-0.16412,1872.6,3950.9,-55.703,-375.73,-9.1004,-19.061
493.0000000000,-0.16406,-686.14,-1835.5,-85.641,-470.30,-9.0975,-18.666
494.0000000000,-0.16410,1870.2,3948.4,-55.698,-375.85,-9.1004,-18.848
495.0000000000,-0.16426,1866.9,3945.0,-55.702,-376.37,-9.1061,-19.068
496.0000000000,-0.16413,-690.95,-1840.6,-85.636,-470.54,-9.1012,-18.697
497.0000000000,-0.16403,-689.05,-1838.6,-85.626,-470.09,-9.0979,-18.675
498.0000000000,-0.16421,1867.5,3945.5,-55.685,-376.01,-9.1051,-19.094
499.0000000000,-0.16416,1864.3,3942.4,-55.690,-376.38,-9.1034,-18.804
500.0000000000,-0.16404,-693.25,-1843.0,-85.624,-470.50,-9.0986,-18.675
501.0000000000,-0.16395,-691.16,-1840.8,-85.613,-470.03,-9.0954,-18.648
502.0000000000,-0.16388,-689.50,-1839.0,-85.606,-469.90,-9.0930,-18.632
503.0000000000,-0.16384,-688.08,-1837.5,-85.600,-469.80,-9.0913,-18.621
504.0000000000,-0.16381,-686.80,-1836.1,-85.593,-469.72,-9.0901,-18.613
505.0000000000,-0.16379,-685.64,-1834.9,-85.586,-469.66,-9.0891,-18.607
506.0000000000,-0.16377,-684.56,-1833.7,-85.580,-469.62,-9.0884,-18.602
507.0000000000,-0.16375,-683.54,-1832.6,-85.573,-469.57,-9.0878,-18.598
508.0000000000,-0.16384,1872.4,3951.0,-55.633,-375.46,-9.0919,-18.775
509.0000000000,-0.16381,-686.07,-1835.2,-85.571,-470.01,-9.0902,-18.630
510.0000000000,-0.16404,1870.5,3948.9,-55.628,-375.68,-9.0989,-19.055
511.0000000000,-0.16568,1867.3,3945.7,-55.631,-377.42,-9.1559,-21.646
512.0000000000,-0.16532,1864.7,3942.9,-55.632,-377.67,-9.1444,-19.304
513.0000000000,-0.16475,-692.77,-1842.2,-85.566,-471.55,-9.1271,-18.916
514.0000000000,-0.16437,-690.66,-1839.9,-85.557,-470.82,-9.1142,-18.813
515.0000000000,-0.16412,-688.91,-1838.0,-85.551,-470.47,-9.1050,-18.752
516.0000000000,-0.16397,-687.45,-1836.4,-85.545,-470.21,-9.0988,-18.710
517.0000000000,-0.16387,-686.10,-1834.9,-85.540,-470.02,-9.0946,-18.680
518.0000000000,-0.16380,-684.87,-1833.6,-85.534,-469.86,-9.0916,-18.658
519.0000000000,-0.16376,-683.73,-1832.4,-85.529,-469.75,-9.0896,-18.642
520.0000000000,-0.16372,-682.68,-1831.3,-85.522,-469.65,-9.0881,-18.629
521.0000000000,-0.16370,-681.70,-1830.2,-85.517,-469.58,-9.0870,-18.620
522.0000000000,-0.16368,-680.76,-1829.1,-85.511,-469.52,-9.0862,-18.612
523.0000000000,-0.16366,-679.84,-1828.2,-85.505,-469.47,-9.0855,-18.606
524.0000000000,-0.16365,-678.95,-1827.2,-85.500,-469.43,-9.0850,-18.602
525.0000000000,-0.16366,1876.9,3956.3,-55.560,-375.25,-9.0864,-18.642
526.0000000000,-0.16366,1873.3,3952.6,-55.565,-375.63,-9.0868,-18.635
527.0000000000,-0.16365,-684.60,-1833.1,-85.499,-469.84,-9.0853,-18.603
528.0000000000,-0.16368,1872.3,3951.4,-55.556,-375.33,-9.0875,-18.693
529.0000000000,-0.16401,1869.3,3948.3,-55.560,-375.94,-9.0989,-19.215
530.0000000000,-0.16456,1866.8,3945.7,-55.561,-376.52,-9.1181,-19.822
531.0000000000,-0.16430,-690.35,-1839.2,-85.494,-470.70,-9.1092,-18.843
532.0000000000,-0.16404,-687.97,-1836.7,-85.484,-470.14,-9.1013,-18.732
533.0000000000,-0.16387,-686.08,-1834.7,-85.477,-469.91,-9.0952,-18.689
534.0000000000,-0.16376,-684.48,-1833.0,-85.471,-469.73,-9.0910,-18.661
535.0000000000,-0.16368,-683.07,-1831.4,-85.465,-469.60,-9.0880,-18.642
536.0000000000,-0.16744,1873.2,3952.5,-55.526,-378.38,-9.2177,-25.150
537.0000000000,-0.16816,1869.4,3949.0,-55.533,-380.35,-9.2438,-22.410
538.0000000000,-0.16727,1866.0,3946.1,-55.541,-380.41,-9.2201,-20.540
539.0000000000,-0.16600,-691.81,-1839.1,-85.483,-473.78,-9.1792,-19.395
540.0000000000,-0.16516,1865.1,3945.7,-55.547,-378.40,-9.1510,-19.198
541.0000000000,-0.16600,1862.2,3942.9,-55.557,-379.14,-9.1777,-21.384
542.0000000000,-0.16534,-695.26,-1842.0,-85.495,-472.93,-9.1523,-19.282
543.0000000000,-0.16473,-693.07,-1839.5,-85.489,-471.93,-9.1317,-19.038
544.0000000000,-0.16436,1863.6,3945.2,-55.552,-377.19,-9.1184,-18.953
545.0000000000,-0.16410,-694.25,-1840.1,-85.493,-471.29,-9.1071,-18.846
546.0000000000,-0.16394,-692.26,-1837.9,-85.486,-470.62,-9.0999,-18.786
547.0000000000,-0.16383,-690.61,-1836.0,-85.483,-470.32,-9.0950,-18.742
548.0000000000,-0.16375,-689.17,-1834.3,-85.479,-470.10,-9.0915,-18.710
549.0000000000,-0.16370,-687.87,-1832.8,-85.476,-469.93,-9.0892,-18.691
550.0000000000,-0.16366,-686.76,-1831.3,-85.471,-469.80,-9.0874,-18.667
551.0000000000,-0.16363,-685.81,-1830.0,-85.467,-469.70,-9.0861,-18.652
552.0000000000,-0.16361,-684.87,-1828.8,-85.463,-469.61,-9.0851,-18.640
553.0000000000,-0.16359,-683.99,-1827.6,-85.458,-469.54,-9.0843,-18.631
554.0000000000,-0.16358,-683.16,-1826.4,-85.452,-469.49,-9.0836,-18.624
555.0000000000,-0.16357,-682.29,-1825.3,-85.447,-469.44,-9.0831,-18.618
556.0000000000,-0.16357,1873.5,3958.3,-55.507,-375.25,-9.0843,-18.644
557.0000000000,-0.16358,1869.9,3954.7,-55.512,-375.63,-9.0848,-18.652
558.0000000000,-0.16386,1867.0,3951.7,-55.514,-375.90,-9.0944,-19.113
559.0000000000,-0.16378,-690.59,-1833.5,-85.449,-470.10,-9.0909,-18.691
560.0000000000,-0.16369,-688.52,-1831.2,-85.439,-469.66,-9.0881,-18.652
561.0000000000,-0.16362,-686.90,-1829.4,-85.433,-469.54,-9.0858,-18.636
562.0000000000,-0.16396,1869.5,3954.7,-55.494,-375.60,-9.0982,-19.275
563.0000000000,-0.16431,1866.3,3951.6,-55.499,-376.33,-9.1102,-19.503
564.0000000000,-0.16442,1863.7,3948.9,-55.501,-376.61,-9.1149,-19.375
565.0000000000,-0.16414,-693.59,-1836.1,-85.436,-470.67,-9.1051,-18.812
566.0000000000,-0.16391,-691.20,-1833.6,-85.426,-470.09,-9.0975,-18.736
567.0000000000,-0.16376,-689.29,-1831.6,-85.421,-469.87,-9.0920,-18.698
568.0000000000,-0.16366,-687.70,-1829.9,-85.416,-469.70,-9.0882,-18.672
569.0000000000,-0.16360,-686.33,-1828.3,-85.411,-469.57,-9.0856,-18.654
570.0000000000,-0.16356,-685.04,-1826.9,-85.407,-469.47,-9.0837,-18.640
571.0000000000,-0.16369,1871.2,3956.9,-55.469,-375.35,-9.0889,-18.906
572.0000000000,-0.16363,-687.08,-1829.0,-85.409,-469.86,-9.0860,-18.667
573.0000000000,-0.16357,-685.34,-1827.2,-85.401,-469.46,-9.0840,-18.641
574.0000000000,-0.16353,-683.91,-1825.7,-85.396,-469.36,-9.0824,-18.629
575.0000000000,-0.16349,-682.61,-1824.3,-85.392,-469.29,-9.0811,-18.620
576.0000000000,-0.16348,-681.41,-1823.1,-85.389,-469.23,-9.0802,-18.614
577.0000000000,-0.16347,-680.29,-1821.9,-85.385,-469.19,-9.0796,-18.609
578.0000000000,-0.16346,-679.24,-1820.8,-85.382,-469.15,-9.0791,-18.607
579.0000000000,-0.16413,1876.8,3962.8,-55.444,-375.50,-9.1029,-19.762
580.0000000000,-0.16574,1873.3,3959.2,-55.451,-377.34,-9.1585,-21.811
581.0000000000,-0.16516,-684.49,-1826.3,-85.387,-471.62,-9.1392,-19.185
582.0000000000,-0.16455,-682.75,-1824.5,-85.379,-470.88,-9.1211,-18.937
583.0000000000,-0.16415,-681.31,-1822.9,-85.376,-470.45,-9.1074,-18.836
584.0000000000,-0.16391,-680.05,-1821.5,-85.372,-470.11,-9.0978,-18.772
585.0000000000,-0.16376,-678.84,-1820.2,-85.369,-469.85,-9.0914,-18.728
586.0000000000,-0.16366,-677.74,-1819.0,-85.365,-469.65,-9.0871,-18.696
587.0000000000,-0.16359,-676.71,-1818.0,-85.360,-469.50,-9.0841,-18.672
588.0000000000,-0.16354,-675.75,-1817.0,-85.355,-469.38,-9.0820,-18.655
589.0000000000,-0.16370,1880.2,3966.5,-55.417,-375.27,-9.0879,-18.954
590.0000000000,-0.16406,1876.7,3962.9,-55.423,-375.95,-9.1005,-19.414
591.0000000000,-0.16390,-681.18,-1822.7,-85.357,-470.13,-9.0943,-18.769
592.0000000000,-0.16373,-679.22,-1820.8,-85.347,-469.63,-9.0892,-18.702
593.0000000000,-0.16363,-677.61,-1819.3,-85.341,-469.46,-9.0854,-18.672
594.0000000000,-0.16366,1878.8,3964.7,-55.401,-375.25,-9.0872,-18.837
595.0000000000,-0.16413,1875.6,3961.3,-55.406,-375.98,-9.1033,-19.594
596.0000000000,-0.16462,1873.0,3958.5,-55.408,-376.54,-9.1203,-19.938
597.0000000000,-0.16429,-684.27,-1826.6,-85.343,-470.66,-9.1088,-18.902
598.0000000000,-0.16397,-681.93,-1824.2,-85.333,-470.04,-9.0990,-18.783
599.0000000000,-0.16377,-680.17,-1822.4,-85.328,-469.76,-9.0918,-18.730
600.0000000000,-0.16365,-678.67,-1820.7,-85.322,-469.55,-9.0868,-18.695
601.0000000000,-0.16356,-677.29,-1819.2,-85.317,-469.39,-9.0833,-18.671
602.0000000000,-0.16351,-676.03,-1817.9,-85.311,-469.26,-9.0809,-18.653
603.0000000000,-0.16347,-674.82,-1816.6,-85.305,-469.17,-9.0792,-18.639
604.0000000000,-0.16344,-673.69,-1815.4,-85.300,-469.09,-9.0780,-18.629
605.0000000000,-0.16344,-672.61,-1814.3,-85.294,-469.03,-9.0775,-18.645
606.0000000000,-0.16342,-671.57,-1813.3,-85.289,-468.98,-9.0767,-18.619
607.0000000000,-0.16348,1884.4,3970.3,-55.350,-374.84,-9.0798,-18.753
608.0000000000,-0.16348,1880.9,3966.7,-55.354,-375.22,-9.0798,-18.670
609.0000000000,-0.16344,-676.88,-1818.9,-85.290,-469.41,-9.0777,-18.625
610.0000000000,-0.16341,-674.92,-1817.0,-85.280,-469.01,-9.0766,-18.615
611.0000000000,-0.16339,-673.35,-1815.4,-85.273,-468.93,-9.0757,-18.609
612.0000000000,-0.16338,-671.98,-1814.0,-85.267,-468.88,-9.0753,-18.622
613.0000000000,-0.16391,1884.2,3969.8,-55.328,-375.11,-9.0942,-19.527
614.0000000000,-0.16393,1881.0,3966.4,-55.333,-375.64,-9.0953,-19.009
615.0000000000,-0.16374,-676.72,-1819.0,-85.268,-469.78,-9.0889,-18.728
616.0000000000,-0.16399,1880.3,3965.6,-55.325,-375.45,-9.0988,-19.364
617.0000000000,-0.16381,-677.44,-1819.9,-85.263,-469.89,-9.0916,-18.767
618.0000000000,-0.16363,-675.37,-1817.8,-85.253,-469.39,-9.0859,-18.700
619.0000000000,-0.16352,-673.69,-1816.0,-85.247,-469.21,-9.0817,-18.669
620.0000000000,-0.16346,-672.22,-1814.5,-85.241,-469.08,-9.0792,-18.672
621.0000000000,-0.16357,1884.1,3969.4,-55.302,-374.94,-9.0835,-18.907
622.0000000000,-0.16362,1880.9,3966.1,-55.307,-375.37,-9.0852,-18.882
623.0000000000,-0.16354,-676.78,-1819.2,-85.242,-469.53,-9.0815,-18.696
624.0000000000,-0.16345,-674.65,-1817.1,-85.232,-469.08,-9.0787,-18.651
625.0000000000,-0.16349,1882.1,3967.2,-55.293,-374.86,-9.0806,-18.792
626.0000000000,-0.16343,-675.84,-1818.4,-85.231,-469.33,-9.0776,-18.653
627.0000000000,-0.16432,1881.1,3966.2,-55.288,-375.51,-9.1090,-20.240
628.0000000000,-0.16416,1878.4,3963.3,-55.292,-375.97,-9.1038,-19.019
629.0000000000,-0.16432,1876.1,3960.9,-55.294,-376.21,-9.1109,-19.568
630.0000000000,-0.16428,1874.0,3958.7,-55.294,-376.30,-9.1100,-19.316
631.0000000000,-0.16396,-682.91,-1826.0,-85.230,-470.26,-9.0985,-18.831
632.0000000000,-0.16372,-680.26,-1823.2,-85.220,-469.63,-9.0899,-18.752
633.0000000000,-0.16357,-678.16,-1821.0,-85.215,-469.37,-9.0842,-18.725
634.0000000000,-0.16349,1878.6,3963.5,-55.275,-375.03,-9.0818,-18.724
635.0000000000,-0.16547,1875.8,3960.6,-55.281,-376.92,-9.1494,-22.178
636.0000000000,-0.16532,1873.5,3958.1,-55.283,-377.35,-9.1447,-19.827
637.0000000000,-0.16464,-683.74,-1826.7,-85.220,-471.21,-9.1237,-19.044
638.0000000000,-0.16415,-681.30,-1824.1,-85.213,-470.38,-9.1072,-18.896
639.0000000000,-0.16383,-679.30,-1822.0,-85.209,-469.94,-9.0955,-18.814
640.0000000000,-0.16364,-677.60,-1820.2,-85.206,-469.62,-9.0877,-18.758
641.0000000000,-0.16351,-676.08,-1818.6,-85.205,-469.38,-9.0823,-18.718
642.0000000000,-0.16343,-674.69,-1817.1,-85.201,-469.19,-9.0787,-18.689
643.0000000000,-0.16338,-673.37,-1815.7,-85.197,-469.04,-9.0761,-18.667
644.0000000000,-0.16334,-672.07,-1814.3,-85.194,-468.93,-9.0743,-18.650
645.0000000000,-0.16331,-670.86,-1813.1,-85.189,-468.83,-9.0730,-18.638
646.0000000000,-0.16329,-669.73,-1811.9,-85.185,-468.76,-9.0720,-18.628
647.0000000000,-0.16327,-668.61,-1810.7,-85.180,-468.70,-9.0713,-18.620
648.0000000000,-0.16326,-667.54,-1809.6,-85.175,-468.65,-9.0707,-18.614
649.0000000000,-0.16410,1888.5,3974.0,-55.236,-375.13,-9.1005,-20.066
650.0000000000,-0.16390,-669.90,-1812.1,-85.176,-469.74,-9.0932,-18.839
651.0000000000,-0.16366,-668.25,-1810.5,-85.168,-469.26,-9.0862,-18.732
652.0000000000,-0.16350,-666.89,-1809.2,-85.163,-469.07,-9.0807,-18.690
653.0000000000,-0.16340,-665.70,-1808.0,-85.159,-468.92,-9.0769,-18.665
654.0000000000,-0.16334,-664.64,-1806.8,-85.154,-468.80,-9.0743,-18.647
655.0000000000,-0.16329,-663.67,-1805.8,-85.149,-468.71,-9.0724,-18.633
656.0000000000,-0.16326,-662.75,-1804.8,-85.144,-468.64,-9.0711,-18.624
657.0000000000,-0.16324,-661.84,-1803.8,-85.139,-468.58,-9.0701,-18.616
658.0000000000,-0.16323,-660.97,-1802.9,-85.134,-468.53,-9.0694,-18.611
659.0000000000,-0.16325,1894.9,3980.6,-55.195,-374.36,-9.0711,-18.667
660.0000000000,-0.16339,1891.3,3976.9,-55.200,-374.85,-9.0761,-18.889
661.0000000000,-0.16383,1888.3,3973.7,-55.202,-375.29,-9.0912,-19.479
662.0000000000,-0.16366,-669.19,-1811.5,-85.139,-469.49,-9.0850,-18.760
663.0000000000,-0.16349,-667.06,-1809.4,-85.130,-469.00,-9.0798,-18.690
664.0000000000,-0.16337,-665.38,-1807.7,-85.125,-468.82,-9.0757,-18.661
665.0000000000,-0.16330,-663.95,-1806.1,-85.120,-468.70,-9.0729,-18.642
666.0000000000,-0.16325,-662.69,-1804.8,-85.116,-468.60,-9.0709,-18.629
667.0000000000,-0.16322,-661.53,-1803.5,-85.110,-468.52,-9.0695,-18.619
668.0000000000,-0.16320,-660.45,-1802.4,-85.105,-468.46,-9.0685,-18.612
669.0000000000,-0.16318,-659.42,-1801.3,-85.100,-468.41,-9.0677,-18.607
670.0000000000,-0.16317,-658.43,-1800.3,-85.095,-468.37,-9.0671,-18.602
671.0000000000,-0.16316,-657.48,-1799.3,-85.090,-468.34,-9.0667,-18.599
672.0000000000,-0.16315,-656.57,-1798.3,-85.085,-468.31,-9.0663,-18.596
673.0000000000,-0.16314,-655.68,-1797.4,-85.080,-468.28,-9.0660,-18.594
674.0000000000,-0.16599,1900.2,3986.0,-55.141,-376.38,-9.1647,-23.483
675.0000000000,-0.16693,1896.6,3982.2,-55.147,-378.30,-9.1982,-22.081
676.0000000000,-0.16585,1893.1,3978.8,-55.151,-378.15,-9.1664,-19.546
677.0000000000,-0.16492,1890.1,3976.0,-55.156,-377.52,-9.1378,-19.207
678.0000000000,-0.16429,-667.42,-1809.1,-85.096,-471.06,-9.1147,-18.996
679.0000000000,-0.16389,-665.32,-1806.9,-85.090,-470.15,-9.0991,-18.888
680.0000000000,-0.16365,-663.64,-1805.1,-85.089,-469.70,-9.0887,-18.815
681.0000000000,-0.16349,-662.25,-1803.6,-85.087,-469.37,-9.0817,-18.762
682.0000000000,-0.16339,-660.99,-1802.2,-85.084,-469.11,-9.0770,-18.722
683.0000000000,-0.16332,-659.78,-1800.8,-85.081,-468.92,-9.0737,-18.693
684.0000000000,-0.16327,-658.62,-1799.6,-85.078,-468.77,-9.0714,-18.670
685.0000000000,-0.16324,-657.54,-1798.4,-85.074,-468.65,-9.0698,-18.653
686.0000000000,-0.16321,-656.52,-1797.3,-85.070,-468.56,-9.0685,-18.640
687.0000000000,-0.16319,-655.54,-1796.3,-85.065,-468.48,-9.0676,-18.630
688.0000000000,-0.16318,-654.61,-1795.3,-85.062,-468.42,-9.0669,-18.621
689.0000000000,-0.16316,-653.73,-1794.4,-85.058,-468.37,-9.0663,-18.615
690.0000000000,-0.16316,-652.91,-1793.5,-85.054,-468.33,-9.0659,-18.610
691.0000000000,-0.16315,-652.16,-1792.6,-85.050,-468.29,-9.0655,-18.607
692.0000000000,-0.16340,1903.5,3990.8,-55.112,-374.31,-9.0751,-19.045
693.0000000000,-0.16334,-655.16,-1795.5,-85.052,-468.86,-9.0722,-18.672
694.0000000000,-0.16326,-653.80,-1794.1,-85.044,-468.47,-9.0699,-18.638
695.0000000000,-0.16321,-652.67,-1792.9,-85.039,-468.38,-9.0681,-18.625
696.0000000000,-0.16318,-651.68,-1791.8,-85.034,-468.31,-9.0667,-18.616
697.0000000000,-0.16315,-650.77,-1790.8,-85.029,-468.26,-9.0658,-18.610
698.0000000000,-0.16314,-649.90,-1789.8,-85.024,-468.22,-9.0650,-18.605
699.0000000000,-0.16312,-649.06,-1789.0,-85.020,-468.18,-9.0645,-18.601
700.0000000000,-0.16311,-648.29,-1788.1,-85.015,-468.15,-9.0641,-18.598
701.0000000000,-0.16310,-647.55,-1787.3,-85.010,-468.13,-9.0637,-18.596
702.0000000000,-0.16309,-646.82,-1786.6,-85.005,-468.11,-9.0634,-18.594
703.0000000000,-0.16308,-646.11,-1785.8,-85.000,-468.08,-9.0631,-18.593
704.0000000000,-0.16308,-645.40,-1785.1,-84.996,-468.06,-9.0628,-18.592
705.0000000000,-0.16307,-644.72,-1784.4,-84.991,-468.05,-9.0626,-18.591
706.0000000000,-0.16306,-644.07,-1783.7,-84.987,-468.03,-9.0624,-18.590
707.0000000000,-0.16306,-643.42,-1783.0,-84.982,-468.01,-9.0622,-18.589
708.0000000000,-0.16305,-642.80,-1782.4,-84.977,-468.00,-9.0620,-18.588
709.0000000000,-0.16305,-642.16,-1781.7,-84.972,-467.99,-9.0619,-18.593
710.0000000000,-0.16305,-641.54,-1781.0,-84.968,-467.98,-9.0621,-18.613
711.0000000000,-0.16304,-640.93,-1780.4,-84.963,-467.97,-9.0618,-18.591
712.0000000000,-0.16304,-640.32,-1779.7,-84.959,-467.95,-9.0615,-18.588
713.0000000000,-0.16303,-639.73,-1779.1,-84.955,-467.93,-9.0612,-18.587
714.0000000000,-0.16302,-639.13,-1778.4,-84.951,-467.92,-9.0609,-18.586
715.0000000000,-0.16301,-638.52,-1777.8,-84.947,-467.90,-9.0606,-18.585
716.0000000000,-0.16301,-637.92,-1777.1,-84.942,-467.89,-9.0604,-18.584
717.0000000000,-0.16300,-637.34,-1776.5,-84.938,-467.87,-9.0602,-18.584
718.0000000000,-0.16303,1918.2,4006.6,-55.000,-373.72,-9.0620,-18.634
719.0000000000,-0.16302,-640.58,-1779.9,-84.941,-468.27,-9.0608,-18.591
720.0000000000,-0.16301,-639.36,-1778.6,-84.933,-467.92,-9.0603,-18.587
721.0000000000,-0.16299,-638.38,-1777.6,-84.929,-467.87,-9.0599,-18.585
722.0000000000,-0.16302,1917.5,4005.8,-54.990,-373.70,-9.0615,-18.632
723.0000000000,-0.16304,1913.9,4002.0,-54.997,-374.11,-9.0625,-18.652
724.0000000000,-0.16302,-644.13,-1783.7,-84.934,-468.32,-9.0610,-18.597
725.0000000000,-0.16300,-642.37,-1782.0,-84.925,-467.93,-9.0602,-18.590
726.0000000000,-0.16298,-641.01,-1780.6,-84.921,-467.87,-9.0595,-18.587
727.0000000000,-0.16407,1915.1,4003.2,-54.982,-374.54,-9.0979,-20.474
728.0000000000,-0.16387,1911.8,3999.7,-54.988,-375.05,-9.0914,-18.970
729.0000000000,-0.16355,-646.02,-1785.9,-84.926,-469.11,-9.0813,-18.763
730.0000000000,-0.16339,1910.9,3998.6,-54.983,-374.43,-9.0771,-18.815
731.0000000000,-0.16345,1908.0,3995.6,-54.989,-374.79,-9.0789,-19.048
732.0000000000,-0.16364,1905.6,3993.0,-54.992,-374.97,-9.0850,-19.289
733.0000000000,-0.16382,1903.4,3990.6,-54.994,-375.19,-9.0912,-19.411
734.0000000000,-0.16356,-653.66,-1794.1,-84.930,-469.23,-9.0817,-18.801
735.0000000000,-0.16334,-651.17,-1791.6,-84.921,-468.64,-9.0743,-18.722
736.0000000000,-0.16320,-649.22,-1789.5,-84.916,-468.40,-9.0689,-18.683
737.0000000000,-0.16311,-647.60,-1787.7,-84.912,-468.22,-9.0652,-18.657
738.0000000000,-0.16305,-646.18,-1786.2,-84.907,-468.08,-9.0625,-18.638
739.0000000000,-0.16303,1910.1,3997.8,-54.968,-373.83,-9.0625,-18.667
740.0000000000,-0.16353,1906.9,3994.5,-54.974,-374.58,-9.0796,-19.533
741.0000000000,-0.16344,1904.3,3991.7,-54.976,-374.67,-9.0767,-18.850
742.0000000000,-0.16327,-653.00,-1793.3,-84.913,-468.75,-9.0705,-18.702
743.0000000000,-0.16314,-650.66,-1791.0,-84.904,-468.24,-9.0661,-18.662
744.0000000000,-0.16306,-648.79,-1789.1,-84.898,-468.07,-9.0628,-18.640
745.0000000000,-0.16300,-647.20,-1787.4,-84.893,-467.94,-9.0605,-18.624
746.0000000000,-0.16296,-645.79,-1786.0,-84.887,-467.85,-9.0589,-18.613
747.0000000000,-0.16293,-644.51,-1784.6,-84.881,-467.78,-9.0577,-18.604
748.0000000000,-0.16291,-643.33,-1783.4,-84.876,-467.73,-9.0569,-18.598
749.0000000000,-0.16290,-642.22,-1782.2,-84.870,-467.68,-9.0562,-18.593
750.0000000000,-0.16288,-641.16,-1781.1,-84.864,-467.64,-9.0557,-18.589
751.0000000000,-0.16287,-640.13,-1780.1,-84.858,-467.61,-9.0553,-18.586
752.0000000000,-0.16322,1915.8,4003.5,-54.918,-373.70,-9.0681,-19.189
753.0000000000,-0.16354,1912.4,3999.8,-54.923,-374.44,-9.0795,-19.377
754.0000000000,-0.16337,1909.5,3996.8,-54.924,-374.50,-9.0747,-18.791
755.0000000000,-0.16319,-647.94,-1788.5,-84.858,-468.57,-9.0681,-18.686
756.0000000000,-0.16306,-645.74,-1786.3,-84.849,-468.06,-9.0636,-18.653
757.0000000000,-0.16297,-643.99,-1784.5,-84.842,-467.90,-9.0604,-18.632
758.0000000000,-0.16292,-642.50,-1783.0,-84.837,-467.78,-9.0581,-18.617
759.0000000000,-0.16288,-641.18,-1781.6,-84.831,-467.69,-9.0565,-18.607
760.0000000000,-0.16285,-639.98,-1780.3,-84.825,-467.63,-9.0554,-18.599
761.0000000000,-0.16316,1916.1,4003.3,-54.885,-373.67,-9.0666,-19.145
762.0000000000,-0.16352,1912.7,3999.8,-54.890,-374.41,-9.0792,-19.441
763.0000000000,-0.16332,-644.99,-1785.7,-84.826,-468.60,-9.0721,-18.757
764.0000000000,-0.16313,-642.99,-1783.7,-84.816,-468.10,-9.0662,-18.684
765.0000000000,-0.16303,1913.6,4000.5,-54.876,-373.77,-9.0636,-18.691
766.0000000000,-0.16294,-644.40,-1785.2,-84.815,-468.20,-9.0595,-18.638
767.0000000000,-0.16289,-642.51,-1783.3,-84.805,-467.76,-9.0570,-18.621
768.0000000000,-0.16285,-640.98,-1781.7,-84.799,-467.65,-9.0553,-18.609
769.0000000000,-0.16282,-639.64,-1780.3,-84.794,-467.57,-9.0540,-18.600
770.0000000000,-0.16280,-638.43,-1779.1,-84.788,-467.50,-9.0531,-18.593
771.0000000000,-0.16278,-637.30,-1777.9,-84.783,-467.46,-9.0524,-18.588
772.0000000000,-0.16277,-636.24,-1776.8,-84.777,-467.42,-9.0518,-18.584
773.0000000000,-0.16276,-635.24,-1775.8,-84.772,-467.38,-9.0514,-18.581
774.0000000000,-0.16275,-634.29,-1774.8,-84.767,-467.36,-9.0510,-18.578
775.0000000000,-0.16274,-633.36,-1773.8,-84.762,-467.33,-9.0506,-18.576
776.0000000000,-0.16273,-632.48,-1772.9,-84.756,-467.31,-9.0503,-18.574
777.0000000000,-0.16273,-631.62,-1772.1,-84.751,-467.29,-9.0503,-18.585
778.0000000000,-0.16276,1924.2,4011.3,-54.811,-373.14,-9.0523,-18.636
779.0000000000,-0.16274,-634.40,-1775.0,-84.751,-467.69,-9.0510,-18.583
780.0000000000,-0.16273,-632.96,-1773.6,-84.742,-467.34,-9.0503,-18.577
781.0000000000,-0.16271,-631.79,-1772.4,-84.737,-467.28,-9.0498,-18.574
782.0000000000,-0.16270,-630.77,-1771.4,-84.731,-467.25,-9.0494,-18.572
783.0000000000,-0.16269,-629.82,-1770.4,-84.726,-467.22,-9.0490,-18.571
784.0000000000,-0.16268,-628.93,-1769.5,-84.721,-467.20,-9.0487,-18.569
785.0000000000,-0.16267,-628.08,-1768.6,-84.716,-467.18,-9.0484,-18.568
786.0000000000,-0.16267,-627.27,-1767.7,-84.711,-467.16,-9.0481,-18.567
787.0000000000,-0.16266,-626.48,-1766.9,-84.705,-467.15,-9.0479,-18.567
788.0000000000,-0.16266,-625.71,-1766.1,-84.700,-467.13,-9.0476,-18.566
789.0000000000,-0.16279,1930.0,4017.1,-54.760,-373.06,-9.0531,-18.794
790.0000000000,-0.16279,1926.3,4013.3,-54.766,-373.49,-9.0535,-18.668
791.0000000000,-0.16276,1923.3,4010.0,-54.767,-373.54,-9.0527,-18.624
792.0000000000,-0.16272,-634.36,-1775.4,-84.703,-467.70,-9.0504,-18.590
793.0000000000,-0.16268,-632.34,-1773.3,-84.693,-467.29,-9.0491,-18.581
794.0000000000,-0.16315,1924.2,4010.8,-54.753,-373.44,-9.0659,-19.413
795.0000000000,-0.16302,-633.82,-1774.9,-84.693,-467.99,-9.0609,-18.707
796.0000000000,-0.16288,-631.97,-1773.1,-84.684,-467.55,-9.0565,-18.644
797.0000000000,-0.16294,1924.5,4011.0,-54.744,-373.38,-9.0595,-18.894
798.0000000000,-0.16288,1921.4,4007.8,-54.749,-373.72,-9.0575,-18.712
799.0000000000,-0.16285,1918.8,4005.0,-54.751,-373.74,-9.0567,-18.739
800.0000000000,-0.16277,-638.45,-1780.0,-84.686,-467.85,-9.0529,-18.627
801.0000000000,-0.16271,-636.12,-1777.6,-84.676,-467.39,-9.0504,-18.607
802.0000000000,-0.16267,-634.28,-1775.7,-84.670,-467.27,-9.0486,-18.595
803.0000000000,-0.16264,-632.70,-1774.0,-84.664,-467.18,-9.0473,-18.586
804.0000000000,-0.16261,-631.32,-1772.5,-84.658,-467.12,-9.0463,-18.580
805.0000000000,-0.16260,-630.06,-1771.2,-84.653,-467.07,-9.0456,-18.575
806.0000000000,-0.16259,-628.90,-1770.0,-84.647,-467.03,-9.0451,-18.571
807.0000000000,-0.16268,1927.2,4013.7,-54.706,-372.92,-9.0492,-18.748
808.0000000000,-0.16266,-631.19,-1772.3,-84.645,-467.47,-9.0477,-18.614
809.0000000000,-0.16317,1925.4,4011.8,-54.702,-373.38,-9.0663,-19.522
810.0000000000,-0.16500,1922.3,4008.6,-54.706,-375.35,-9.1296,-22.127
811.0000000000,-0.16552,1919.7,4005.8,-54.707,-376.39,-9.1492,-21.142
812.0000000000,-0.16461,-637.92,-1779.4,-84.644,-470.30,-9.1208,-19.237
813.0000000000,-0.16386,-635.93,-1777.1,-84.636,-469.34,-9.0971,-18.989
814.0000000000,-0.16339,-634.30,-1775.2,-84.632,-468.77,-9.0800,-18.869
815.0000000000,-0.16316,1922.2,4009.0,-54.693,-374.22,-9.0717,-18.908
816.0000000000,-0.16296,-635.91,-1776.7,-84.634,-468.44,-9.0625,-18.753
817.0000000000,-0.16282,-634.09,-1774.8,-84.626,-467.85,-9.0566,-18.704
818.0000000000,-0.16273,-632.56,-1773.3,-84.622,-467.63,-9.0525,-18.670
819.0000000000,-0.16267,-631.20,-1771.8,-84.618,-467.46,-9.0497,-18.646
820.0000000000,-0.16263,-630.00,-1770.5,-84.613,-467.33,-9.0477,-18.627
821.0000000000,-0.16260,-628.87,-1769.3,-84.609,-467.22,-9.0462,-18.612
822.0000000000,-0.16257,-627.81,-1768.2,-84.604,-467.14,-9.0452,-18.601
823.0000000000,-0.16256,-626.80,-1767.1,-84.599,-467.08,-9.0443,-18.593
824.0000000000,-0.16254,-625.83,-1766.0,-84.594,-467.02,-9.0437,-18.586
825.0000000000,-0.16253,-624.95,-1765.0,-84.589,-466.98,-9.0432,-18.581
826.0000000000,-0.16262,1931.0,4018.5,-54.649,-372.86,-9.0472,-18.746
827.0000000000,-0.16259,-627.56,-1767.7,-84.589,-467.40,-9.0454,-18.601
828.0000000000,-0.16259,1928.9,4016.3,-54.645,-372.89,-9.0462,-18.632
829.0000000000,-0.16279,1925.8,4012.9,-54.650,-373.41,-9.0534,-18.987
830.0000000000,-0.16271,-631.90,-1772.5,-84.587,-467.61,-9.0500,-18.645
831.0000000000,-0.16263,-629.86,-1770.4,-84.578,-467.18,-9.0473,-18.611
832.0000000000,-0.16274,1926.7,4013.8,-54.638,-373.04,-9.0518,-18.871
833.0000000000,-0.16354,1923.7,4010.7,-54.644,-374.07,-9.0794,-20.124
834.0000000000,-0.16328,-633.90,-1774.5,-84.581,-468.30,-9.0699,-18.844
835.0000000000,-0.16299,-631.81,-1772.3,-84.572,-467.75,-9.0613,-18.725
836.0000000000,-0.16325,1924.8,4012.0,-54.633,-373.71,-9.0713,-19.453
837.0000000000,-0.16315,1921.8,4009.0,-54.638,-374.05,-9.0674,-18.959
838.0000000000,-0.16360,1919.3,4006.4,-54.640,-374.47,-9.0834,-19.883
839.0000000000,-0.16331,1917.1,4004.1,-54.642,-374.39,-9.0735,-18.891
840.0000000000,-0.16302,-639.93,-1780.5,-84.578,-468.33,-9.0631,-18.753
841.0000000000,-0.16282,-637.43,-1777.8,-84.569,-467.71,-9.0559,-18.699
842.0000000000,-0.16270,-635.46,-1775.7,-84.564,-467.47,-9.0509,-18.664
843.0000000000,-0.16262,-633.78,-1773.8,-84.559,-467.29,-9.0475,-18.639
844.0000000000,-0.16306,1922.7,4010.5,-54.621,-373.39,-9.0631,-19.467
845.0000000000,-0.16292,-635.31,-1775.1,-84.561,-467.89,-9.0570,-18.743
846.0000000000,-0.16276,-633.37,-1773.1,-84.553,-467.41,-9.0519,-18.672
847.0000000000,-0.16348,1923.2,4011.1,-54.613,-373.74,-9.0775,-20.061
848.0000000000,-0.16323,-634.77,-1774.5,-84.553,-468.25,-9.0679,-18.848
849.0000000000,-0.16295,-632.86,-1772.5,-84.544,-467.71,-9.0594,-18.732
850.0000000000,-0.16277,-631.32,-1770.8,-84.538,-467.47,-9.0530,-18.683
851.0000000000,-0.16265,-630.01,-1769.4,-84.534,-467.29,-9.0486,-18.652
852.0000000000,-0.16258,-628.77,-1768.0,-84.530,-467.14,-9.0454,-18.630
853.0000000000,-0.16253,-627.62,-1766.8,-84.525,-467.03,-9.0433,-18.613
854.0000000000,-0.16250,-626.54,-1765.6,-84.521,-466.94,-9.0418,-18.601
855.0000000000,-0.16248,-625.50,-1764.4,-84.516,-466.88,-9.0410,-18.604
856.0000000000,-0.16247,-624.51,-1763.4,-84.512,-466.83,-9.0401,-18.587
857.0000000000,-0.16247,1931.4,4020.2,-54.573,-372.64,-9.0412,-18.615
858.0000000000,-0.16246,-627.05,-1766.0,-84.513,-467.16,-9.0398,-18.582
859.0000000000,-0.16244,-625.52,-1764.4,-84.504,-466.80,-9.0392,-18.576
860.0000000000,-0.16243,-624.25,-1763.1,-84.499,-466.74,-9.0386,-18.572
861.0000000000,-0.16499,1931.9,4020.6,-54.560,-374.59,-9.1273,-22.972
862.0000000000,-0.16631,1928.5,4017.1,-54.565,-376.72,-9.1736,-22.513
863.0000000000,-0.16656,1925.1,4013.9,-54.570,-377.71,-9.1875,-21.854
864.0000000000,-0.16580,1922.0,4011.1,-54.575,-377.61,-9.1654,-20.409
865.0000000000,-0.16495,1919.3,4008.6,-54.582,-377.06,-9.1384,-19.802
866.0000000000,-0.16517,1916.9,4006.3,-54.590,-377.14,-9.1454,-20.993
867.0000000000,-0.16626,1914.7,4004.1,-54.599,-378.07,-9.1817,-22.547
868.0000000000,-0.16519,-642.91,-1780.6,-84.542,-471.72,-9.1439,-19.568
869.0000000000,-0.16425,-640.85,-1778.0,-84.542,-470.48,-9.1130,-19.227
870.0000000000,-0.16363,-639.23,-1775.9,-84.546,-469.66,-9.0903,-19.040
871.0000000000,-0.16408,1917.2,4008.6,-54.615,-375.53,-9.1044,-20.353
872.0000000000,-0.16383,1914.1,4005.8,-54.627,-375.66,-9.0941,-19.365
873.0000000000,-0.16345,1911.5,4003.4,-54.635,-375.30,-9.0810,-19.032
874.0000000000,-0.16363,1908.9,4001.3,-54.642,-375.31,-9.0867,-19.709
875.0000000000,-0.16336,1906.5,3999.4,-54.648,-375.06,-9.0765,-19.004
876.0000000000,-0.16329,1904.3,3997.6,-54.653,-374.90,-9.0740,-19.185
877.0000000000,-0.16305,-652.70,-1786.6,-84.592,-468.79,-9.0643,-18.821
878.0000000000,-0.16287,-650.13,-1783.5,-84.586,-468.13,-9.0574,-18.752
879.0000000000,-0.16490,1906.9,4001.5,-54.650,-375.41,-9.1275,-22.399
880.0000000000,-0.16438,1904.2,3998.9,-54.659,-375.85,-9.1100,-19.335
881.0000000000,-0.16540,1901.5,3996.7,-54.667,-376.81,-9.1484,-21.864
882.0000000000,-0.16459,-655.68,-1787.9,-84.610,-470.70,-9.1204,-19.334
883.0000000000,-0.16386,-653.61,-1785.2,-84.610,-469.72,-9.0968,-19.053
884.0000000000,-0.16338,-651.96,-1783.0,-84.613,-469.11,-9.0797,-18.924
885.0000000000,-0.16308,-650.56,-1781.1,-84.617,-468.65,-9.0679,-18.839
886.0000000000,-0.16290,-649.21,-1779.4,-84.621,-468.30,-9.0601,-18.779
887.0000000000,-0.16279,-647.91,-1777.7,-84.623,-468.04,-9.0548,-18.735
888.0000000000,-0.16271,-646.63,-1776.1,-84.624,-467.84,-9.0512,-18.702
889.0000000000,-0.16266,-645.47,-1774.7,-84.625,-467.67,-9.0486,-18.677
890.0000000000,-0.16263,-644.40,-1773.4,-84.627,-467.55,-9.0469,-18.658
891.0000000000,-0.16261,-643.49,-1772.1,-84.629,-467.46,-9.0457,-18.643
892.0000000000,-0.16259,-642.68,-1770.9,-84.630,-467.38,-9.0448,-18.632
893.0000000000,-0.16258,-641.80,-1769.8,-84.628,-467.32,-9.0441,-18.623
894.0000000000,-0.16275,1914.1,4013.8,-54.693,-373.25,-9.0507,-18.918
895.0000000000,-0.16413,1910.6,4010.3,-54.702,-374.76,-9.0980,-21.092
896.0000000000,-0.16392,1907.6,4007.3,-54.708,-375.04,-9.0918,-19.293
897.0000000000,-0.16414,1905.1,4004.6,-54.713,-375.38,-9.1018,-20.040
898.0000000000,-0.16395,1902.7,4002.2,-54.718,-375.40,-9.0961,-19.463
899.0000000000,-0.16354,1900.5,4000.0,-54.723,-375.13,-9.0827,-18.986
900.0000000000,-0.16323,1898.5,3997.9,-54.729,-374.82,-9.0717,-18.854
901.0000000000,-0.16367,1896.6,3996.0,-54.734,-375.07,-9.0861,-19.898
902.0000000000,-0.16345,1894.8,3994.2,-54.739,-374.96,-9.0780,-19.026
903.0000000000,-0.16317,-661.74,-1790.0,-84.677,-468.87,-9.0674,-18.813
904.0000000000,-0.16313,1896.2,3995.5,-54.736,-374.19,-9.0667,-19.036
905.0000000000,-0.16297,-660.97,-1789.3,-84.678,-468.50,-9.0599,-18.772
906.0000000000,-0.16285,-658.39,-1786.6,-84.673,-467.96,-9.0550,-18.712
907.0000000000,-0.16276,-656.28,-1784.3,-84.671,-467.76,-9.0514,-18.682
908.0000000000,-0.16355,1900.6,4000.2,-54.735,-374.13,-9.0790,-20.111
909.0000000000,-0.16410,1897.8,3997.3,-54.744,-375.11,-9.0977,-20.194
910.0000000000,-0.16371,1895.6,3995.0,-54.749,-375.08,-9.0860,-19.045
911.0000000000,-0.16333,-661.43,-1789.7,-84.688,-468.98,-9.0730,-18.850
912.0000000000,-0.16327,1896.1,3995.5,-54.749,-374.31,-9.0716,-19.117
913.0000000000,-0.16307,-661.19,-1789.4,-84.692,-468.60,-9.0629,-18.783
914.0000000000,-0.16291,-658.68,-1786.8,-84.685,-468.03,-9.0569,-18.726
915.0000000000,-0.16281,-656.62,-1784.7,-84.682,-467.82,-9.0528,-18.694
916.0000000000,-0.16274,-654.77,-1782.8,-84.679,-467.66,-9.0498,-18.670
917.0000000000,-0.16270,-653.11,-1781.2,-84.677,-467.54,-9.0478,-18.653
918.0000000000,-0.16267,-651.56,-1779.7,-84.676,-467.45,-9.0466,-18.650
919.0000000000,-0.16352,1904.8,4004.3,-54.739,-373.91,-9.0763,-20.114
920.0000000000,-0.16331,-653.21,-1781.6,-84.681,-468.49,-9.0685,-18.861
921.0000000000,-0.16306,-651.27,-1779.7,-84.674,-468.00,-9.0611,-18.749
922.0000000000,-0.16289,-649.60,-1778.2,-84.669,-467.79,-9.0554,-18.704
923.0000000000,-0.16278,-648.11,-1776.8,-84.664,-467.62,-9.0514,-18.676
924.0000000000,-0.16271,-646.78,-1775.5,-84.659,-467.50,-9.0486,-18.656
925.0000000000,-0.16266,-645.57,-1774.4,-84.655,-467.40,-9.0467,-18.641
926.0000000000,-0.16263,-644.39,-1773.3,-84.650,-467.32,-9.0454,-18.631
927.0000000000,-0.16260,-643.24,-1772.2,-84.646,-467.26,-9.0444,-18.622
928.0000000000,-0.16259,-642.17,-1771.2,-84.642,-467.21,-9.0437,-18.616
929.0000000000,-0.16257,-641.14,-1770.2,-84.638,-467.17,-9.0431,-18.611
930.0000000000,-0.16256,-640.14,-1769.3,-84.633,-467.14,-9.0427,-18.607
931.0000000000,-0.16255,-639.17,-1768.3,-84.628,-467.11,-9.0423,-18.604
932.0000000000,-0.16254,-638.24,-1767.4,-84.623,-467.09,-9.0420,-18.602
933.0000000000,-0.16253,-637.33,-1766.5,-84.618,-467.07,-9.0417,-18.600
934.0000000000,-0.16252,-636.42,-1765.7,-84.613,-467.05,-9.0415,-18.598
935.0000000000,-0.16251,-635.50,-1764.8,-84.608,-467.03,-9.0412,-18.597
936.0000000000,-0.16250,-634.60,-1764.0,-84.604,-467.01,-9.0410,-18.595
937.0000000000,-0.16250,-633.71,-1763.2,-84.600,-466.99,-9.0408,-18.594
938.0000000000,-0.16249,-632.84,-1762.4,-84.595,-466.98,-9.0406,-18.593
939.0000000000,-0.16248,-631.98,-1761.6,-84.590,-466.96,-9.0404,-18.592
940.0000000000,-0.16247,-631.12,-1760.9,-84.585,-466.95,-9.0401,-18.592
941.0000000000,-0.16247,-630.25,-1760.2,-84.581,-466.94,-9.0399,-18.591
942.0000000000,-0.16246,-629.39,-1759.5,-84.576,-466.92,-9.0397,-18.590
943.0000000000,-0.16269,1926.5,4023.7,-54.637,-372.94,-9.0488,-19.001
944.0000000000,-0.16288,1922.9,4019.7,-54.644,-373.54,-9.0554,-19.074
945.0000000000,-0.16276,-635.06,-1766.1,-84.581,-467.75,-9.0508,-18.693
946.0000000000,-0.16264,-633.23,-1764.5,-84.573,-467.31,-9.0471,-18.652
947.0000000000,-0.16256,-631.76,-1763.1,-84.569,-467.18,-9.0444,-18.633
948.0000000000,-0.16251,-630.50,-1761.9,-84.565,-467.09,-9.0424,-18.620
949.0000000000,-0.16248,-629.35,-1760.9,-84.562,-467.02,-9.0410,-18.612
950.0000000000,-0.16246,-628.29,-1759.9,-84.557,-466.97,-9.0400,-18.605
951.0000000000,-0.16244,-627.30,-1759.0,-84.552,-466.93,-9.0393,-18.601
952.0000000000,-0.16243,-626.35,-1758.1,-84.547,-466.89,-9.0387,-18.597
953.0000000000,-0.16242,-625.44,-1757.3,-84.542,-466.86,-9.0383,-18.594
954.0000000000,-0.16241,-624.57,-1756.5,-84.536,-466.84,-9.0379,-18.591
955.0000000000,-0.16264,1931.3,4026.7,-54.596,-372.85,-9.0469,-19.005
956.0000000000,-0.16276,1927.7,4022.9,-54.601,-373.39,-9.0514,-18.968
957.0000000000,-0.16302,1924.7,4019.6,-54.603,-373.72,-9.0607,-19.303
958.0000000000,-0.16337,1922.1,4016.7,-54.604,-374.14,-9.0732,-19.646
959.0000000000,-0.16308,-635.18,-1768.4,-84.539,-468.25,-9.0633,-18.825
960.0000000000,-0.16283,-632.87,-1766.1,-84.529,-467.68,-9.0553,-18.733
961.0000000000,-0.16267,-631.06,-1764.3,-84.523,-467.43,-9.0493,-18.690
962.0000000000,-0.16330,1925.4,4019.8,-54.582,-373.68,-9.0711,-19.914
963.0000000000,-0.16340,1922.3,4016.5,-54.587,-374.27,-9.0742,-19.393
964.0000000000,-0.16309,-635.20,-1768.8,-84.523,-468.32,-9.0634,-18.828
965.0000000000,-0.16284,-633.01,-1766.7,-84.513,-467.73,-9.0551,-18.744
966.0000000000,-0.16269,-631.29,-1765.0,-84.507,-467.47,-9.0491,-18.700
967.0000000000,-0.16258,-629.87,-1763.5,-84.501,-467.28,-9.0449,-18.671
968.0000000000,-0.16266,1926.4,4020.4,-54.562,-373.08,-9.0477,-18.889
969.0000000000,-0.16276,1923.2,4017.0,-54.567,-373.53,-9.0510,-18.975
970.0000000000,-0.16265,-634.48,-1768.4,-84.502,-467.67,-9.0464,-18.693
971.0000000000,-0.16255,-632.34,-1766.3,-84.493,-467.19,-9.0430,-18.655
972.0000000000,-0.16249,-630.60,-1764.6,-84.486,-467.05,-9.0405,-18.636
973.0000000000,-0.16255,1925.9,4019.5,-54.546,-372.86,-9.0430,-18.786
974.0000000000,-0.16251,-632.21,-1766.3,-84.485,-467.35,-9.0402,-18.640
975.0000000000,-0.16247,-630.34,-1764.5,-84.476,-466.95,-9.0385,-18.621
976.0000000000,-0.16244,-628.81,-1762.9,-84.470,-466.85,-9.0371,-18.610
977.0000000000,-0.16242,-627.47,-1761.5,-84.465,-466.79,-9.0361,-18.603
978.0000000000,-0.16241,-626.24,-1760.2,-84.459,-466.74,-9.0354,-18.598
979.0000000000,-0.16241,-625.08,-1759.1,-84.454,-466.70,-9.0348,-18.594
980.0000000000,-0.16240,-624.00,-1758.0,-84.449,-466.67,-9.0344,-18.590
981.0000000000,-0.16240,-622.97,-1757.0,-84.443,-466.64,-9.0340,-18.588
982.0000000000,-0.16240,-622.00,-1755.9,-84.437,-466.61,-9.0337,-18.586
983.0000000000,-0.16282,1933.9,4027.6,-54.497,-372.77,-9.0489,-19.311
984.0000000000,-0.16272,-624.53,-1758.6,-84.435,-467.35,-9.0449,-18.702
985.0000000000,-0.16285,1932.0,4025.4,-54.491,-372.98,-9.0508,-19.073
986.0000000000,-0.16272,-626.06,-1760.5,-84.430,-467.45,-9.0455,-18.695
987.0000000000,-0.16260,-624.23,-1758.7,-84.420,-467.00,-9.0415,-18.651
988.0000000000,-0.16253,-622.73,-1757.3,-84.413,-466.86,-9.0385,-18.631
989.0000000000,-0.16248,-621.40,-1756.0,-84.407,-466.77,-9.0364,-18.617
990.0000000000,-0.16244,-620.19,-1754.9,-84.401,-466.69,-9.0349,-18.607
991.0000000000,-0.16241,-619.09,-1753.9,-84.395,-466.63,-9.0338,-18.599
992.0000000000,-0.16239,-618.10,-1752.9,-84.389,-466.58,-9.0330,-18.594
993.0000000000,-0.16238,-617.15,-1751.9,-84.383,-466.55,-9.0324,-18.590
994.0000000000,-0.16236,-616.24,-1751.1,-84.377,-466.51,-9.0319,-18.586
995.0000000000,-0.16235,-615.35,-1750.2,-84.371,-466.48,-9.0315,-18.584
996.0000000000,-0.16234,-614.50,-1749.4,-84.365,-466.46,-9.0312,-18.581
997.0000000000,-0.16233,-613.67,-1748.7,-84.359,-466.44,-9.0308,-18.580
998.0000000000,-0.16232,-612.86,-1747.9,-84.353,-466.42,-9.0306,-18.578
999.0000000000,-0.16232,-612.07,-1747.2,-84.347,-466.40,-9.0303,-18.577
1000.000000000,-0.16248,1945.2,4036.1,-54.407,-372.36,-9.0370,-18.875
1001.000000000,-0.16244,-614.77,-1750.3,-84.345,-466.92,-9.0348,-18.624
1002.000000000,-0.16238,-613.45,-1749.0,-84.335,-466.55,-9.0331,-18.601
1003.000000000,-0.16234,-612.35,-1747.9,-84.328,-466.48,-9.0318,-18.592
1004.000000000,-0.16231,-611.36,-1746.9,-84.322,-466.43,-9.0308,-18.587
1005.000000000,-0.16229,-610.44,-1746.0,-84.316,-466.39,-9.0300,-18.582
1006.000000000,-0.16228,-609.58,-1745.1,-84.309,-466.36,-9.0295,-18.579
1007.000000000,-0.16227,-608.76,-1744.3,-84.303,-466.33,-9.0290,-18.577
1008.000000000,-0.16226,-607.96,-1743.5,-84.297,-466.31,-9.0286,-18.575
1009.000000000,-0.16225,-607.18,-1742.8,-84.291,-466.29,-9.0285,-18.582
1010.000000000,-0.16224,-606.43,-1742.0,-84.285,-466.27,-9.0282,-18.574
1011.000000000,-0.16223,-605.71,-1741.3,-84.279,-466.25,-9.0279,-18.572
1012.000000000,-0.16421,1953.2,4041.9,-54.338,-373.67,-9.0966,-21.978
1013.000000000,-0.16407,1947.3,4038.0,-54.343,-374.49,-9.0926,-19.647
1014.000000000,-0.16344,-611.50,-1747.8,-84.279,-468.46,-9.0740,-18.956
1015.000000000,-0.16299,-609.94,-1746.2,-84.269,-467.72,-9.0594,-18.826
1016.000000000,-0.16271,-608.68,-1744.8,-84.264,-467.35,-9.0490,-18.755
1017.000000000,-0.16253,-607.59,-1743.7,-84.259,-467.07,-9.0419,-18.708
1018.000000000,-0.16242,-606.60,-1742.6,-84.254,-466.86,-9.0371,-18.674
1019.000000000,-0.16234,-605.71,-1741.7,-84.249,-466.69,-9.0338,-18.649
1020.000000000,-0.16229,-604.92,-1740.8,-84.244,-466.57,-9.0316,-18.630
1021.000000000,-0.16226,-604.17,-1739.9,-84.239,-466.47,-9.0300,-18.616
1022.000000000,-0.16223,-603.44,-1739.1,-84.234,-466.40,-9.0288,-18.605
1023.000000000,-0.16221,-602.75,-1738.3,-84.229,-466.34,-9.0279,-18.597
1024.000000000,-0.16220,-602.10,-1737.6,-84.224,-466.29,-9.0272,-18.591
1025.000000000,-0.16231,1957.5,4045.6,-54.285,-372.19,-9.0320,-18.798
1026.000000000,-0.16249,1952.0,4041.7,-54.290,-372.74,-9.0384,-18.991
1027.000000000,-0.16650,1948.2,4038.4,-54.293,-376.07,-9.1764,-25.714
1028.000000000,-0.16730,1944.9,4035.2,-54.297,-377.88,-9.2053,-22.845
1029.000000000,-0.16571,-613.83,-1750.1,-84.238,-471.60,-9.1574,-19.724
1030.000000000,-0.16443,-612.38,-1748.2,-84.235,-470.26,-9.1173,-19.304
1031.000000000,-0.16362,-611.25,-1746.7,-84.238,-469.33,-9.0883,-19.099
1032.000000000,-0.16312,-610.30,-1745.3,-84.241,-468.61,-9.0686,-18.964
1033.000000000,-0.16297,1947.4,4038.6,-54.306,-374.04,-9.0620,-19.145
1034.000000000,-0.16514,1942.9,4035.2,-54.315,-375.96,-9.1345,-22.963
1035.000000000,-0.16443,-615.29,-1750.1,-84.253,-470.09,-9.1089,-19.431
1036.000000000,-0.16365,-613.90,-1748.2,-84.249,-469.13,-9.0851,-19.090
1037.000000000,-0.16314,-612.69,-1746.5,-84.249,-468.50,-9.0672,-18.947
1038.000000000,-0.16282,-611.67,-1745.1,-84.248,-468.00,-9.0547,-18.854
1039.000000000,-0.16262,-610.81,-1743.8,-84.246,-467.62,-9.0462,-18.788
1040.000000000,-0.16250,-610.01,-1742.6,-84.245,-467.34,-9.0405,-18.740
1041.000000000,-0.16251,1947.3,4041.0,-54.309,-373.04,-9.0411,-18.879
1042.000000000,-0.16253,1942.5,4037.4,-54.317,-373.35,-9.0411,-18.863
1043.000000000,-0.16244,-615.78,-1748.1,-84.255,-467.44,-9.0369,-18.699
1044.000000000,-0.16237,-614.26,-1746.1,-84.247,-466.95,-9.0341,-18.666
1045.000000000,-0.16232,-613.02,-1744.4,-84.242,-466.80,-9.0321,-18.647
1046.000000000,-0.16229,-612.00,-1743.0,-84.239,-466.69,-9.0305,-18.632
1047.000000000,-0.16226,-611.09,-1741.8,-84.235,-466.61,-9.0294,-18.622
1048.000000000,-0.16230,1945.9,4041.9,-54.298,-372.43,-9.0314,-18.700
1049.000000000,-0.16245,1941.4,4038.3,-54.304,-372.92,-9.0367,-18.921
1050.000000000,-0.16242,1938.3,4035.3,-54.307,-372.98,-9.0358,-18.714
1051.000000000,-0.16241,1935.6,4032.6,-54.310,-373.01,-9.0357,-18.740
1052.000000000,-0.16234,-621.67,-1752.3,-84.248,-467.13,-9.0326,-18.640
1053.000000000,-0.16229,-619.46,-1749.9,-84.241,-466.69,-9.0306,-18.623
1054.000000000,-0.16225,-617.71,-1748.0,-84.238,-466.58,-9.0292,-18.612
1055.000000000,-0.16222,-616.33,-1746.3,-84.236,-466.51,-9.0281,-18.605
1056.000000000,-0.16220,-615.13,-1744.9,-84.233,-466.46,-9.0273,-18.600
1057.000000000,-0.16219,-614.04,-1743.6,-84.230,-466.42,-9.0267,-18.596
1058.000000000,-0.16217,-613.01,-1742.4,-84.228,-466.38,-9.0262,-18.592
1059.000000000,-0.16217,-612.07,-1741.2,-84.227,-466.35,-9.0258,-18.590
1060.000000000,-0.16224,1944.5,4042.4,-54.291,-372.23,-9.0292,-18.716
1061.000000000,-0.16258,1940.5,4038.8,-54.299,-372.90,-9.0408,-19.218
1062.000000000,-0.16398,1937.6,4035.7,-54.304,-374.17,-9.0887,-21.256
1063.000000000,-0.16360,1935.0,4033.1,-54.309,-374.33,-9.0768,-19.167
1064.000000000,-0.16311,-622.30,-1751.9,-84.247,-468.23,-9.0613,-18.872
1065.000000000,-0.16277,-620.18,-1749.6,-84.240,-467.54,-9.0498,-18.783
1066.000000000,-0.16256,-618.46,-1747.6,-84.236,-467.21,-9.0418,-18.729
1067.000000000,-0.16243,-616.93,-1746.0,-84.232,-466.98,-9.0364,-18.692
1068.000000000,-0.16235,-615.71,-1744.5,-84.227,-466.80,-9.0328,-18.665
1069.000000000,-0.16229,-614.58,-1743.2,-84.222,-466.67,-9.0303,-18.645
1070.000000000,-0.16226,-613.50,-1742.0,-84.218,-466.56,-9.0285,-18.630
1071.000000000,-0.16223,-612.47,-1740.9,-84.214,-466.48,-9.0273,-18.619
1072.000000000,-0.16221,-611.58,-1739.9,-84.210,-466.42,-9.0264,-18.610
1073.000000000,-0.16220,-610.74,-1738.9,-84.205,-466.37,-9.0257,-18.604
1074.000000000,-0.16219,-609.92,-1737.9,-84.201,-466.33,-9.0252,-18.598
1075.000000000,-0.16218,-609.16,-1737.1,-84.196,-466.29,-9.0247,-18.594
1076.000000000,-0.16217,-608.42,-1736.2,-84.191,-466.26,-9.0244,-18.591
1077.000000000,-0.16392,1948.9,4047.1,-54.252,-373.48,-9.0851,-21.592
1078.000000000,-0.16352,-611.07,-1739.2,-84.192,-468.18,-9.0712,-19.066
1079.000000000,-0.16304,-609.89,-1737.7,-84.184,-467.59,-9.0574,-18.850
1080.000000000,-0.16272,-608.93,-1736.5,-84.179,-467.26,-9.0467,-18.768
1081.000000000,-0.16252,-608.10,-1735.5,-84.174,-466.99,-9.0393,-18.718
1082.000000000,-0.16240,-607.24,-1734.5,-84.170,-466.79,-9.0342,-18.683
1083.000000000,-0.16232,-606.42,-1733.5,-84.165,-466.63,-9.0307,-18.658
1084.000000000,-0.16227,-605.64,-1732.6,-84.161,-466.51,-9.0284,-18.640
1085.000000000,-0.16223,-604.88,-1731.8,-84.156,-466.42,-9.0268,-18.626
1086.000000000,-0.16221,-604.18,-1731.0,-84.152,-466.35,-9.0256,-18.615
1087.000000000,-0.16219,-603.51,-1730.2,-84.148,-466.29,-9.0247,-18.607
1088.000000000,-0.16218,-602.84,-1729.4,-84.144,-466.24,-9.0241,-18.600
1089.000000000,-0.16217,-602.18,-1728.7,-84.140,-466.21,-9.0236,-18.595
1090.000000000,-0.16216,-601.52,-1728.0,-84.136,-466.17,-9.0232,-18.592
1091.000000000,-0.16364,1957.9,4055.2,-54.197,-373.17,-9.0747,-21.135
1092.000000000,-0.16361,1952.2,4051.3,-54.204,-373.94,-9.0742,-19.516
1093.000000000,-0.16312,-607.17,-1734.6,-84.141,-467.96,-9.0594,-18.893
1094.000000000,-0.16276,-605.62,-1732.9,-84.133,-467.30,-9.0479,-18.786
1095.000000000,-0.16254,-604.44,-1731.6,-84.129,-467.00,-9.0396,-18.729
1096.000000000,-0.16240,-603.49,-1730.5,-84.124,-466.77,-9.0340,-18.690
1097.000000000,-0.16233,1955.6,4053.1,-54.187,-372.45,-9.0318,-18.697
1098.000000000,-0.16253,1950.5,4049.4,-54.193,-372.94,-9.0386,-19.113
1099.000000000,-0.16243,-608.53,-1736.2,-84.131,-467.09,-9.0339,-18.706
1100.000000000,-0.16232,-606.89,-1734.4,-84.123,-466.61,-9.0302,-18.661
1101.000000000,-0.16225,-605.54,-1732.8,-84.118,-466.46,-9.0275,-18.639
1102.000000000,-0.16220,-604.39,-1731.5,-84.115,-466.35,-9.0255,-18.624
1103.000000000,-0.16217,-603.36,-1730.3,-84.111,-466.27,-9.0241,-18.613
1104.000000000,-0.16214,-602.43,-1729.2,-84.107,-466.20,-9.0231,-18.604
1105.000000000,-0.16212,-601.57,-1728.2,-84.103,-466.15,-9.0224,-18.598
1106.000000000,-0.16211,-600.77,-1727.3,-84.099,-466.11,-9.0218,-18.593
1107.000000000,-0.16210,-600.01,-1726.4,-84.095,-466.07,-9.0214,-18.589
1108.000000000,-0.16209,-599.29,-1725.5,-84.091,-466.04,-9.0210,-18.586
1109.000000000,-0.16208,-598.61,-1724.7,-84.086,-466.02,-9.0207,-18.584
1110.000000000,-0.16207,-597.97,-1723.9,-84.081,-466.00,-9.0204,-18.582
1111.000000000,-0.16206,-597.35,-1723.2,-84.077,-465.98,-9.0201,-18.580
1112.000000000,-0.16206,-596.75,-1722.5,-84.072,-465.96,-9.0199,-18.579
1113.000000000,-0.16205,-596.17,-1721.7,-84.067,-465.94,-9.0197,-18.578
1114.000000000,-0.16204,-595.60,-1721.0,-84.063,-465.93,-9.0195,-18.577
1115.000000000,-0.16204,-595.04,-1720.4,-84.058,-465.91,-9.0193,-18.576
1116.000000000,-0.16203,-594.49,-1719.7,-84.053,-465.90,-9.0191,-18.575
1117.000000000,-0.16203,-593.94,-1719.1,-84.048,-465.88,-9.0189,-18.574
1118.000000000,-0.16202,-593.41,-1718.4,-84.043,-465.87,-9.0187,-18.573
1119.000000000,-0.16201,-592.88,-1717.8,-84.038,-465.86,-9.0186,-18.573
1120.000000000,-0.16201,-592.37,-1717.2,-84.033,-465.84,-9.0184,-18.572
1121.000000000,-0.16200,-591.87,-1716.6,-84.027,-465.83,-9.0182,-18.572
1122.000000000,-0.16290,1967.7,4066.5,-54.088,-372.38,-9.0501,-20.125
1123.000000000,-0.16269,-595.12,-1720.0,-84.027,-467.02,-9.0425,-18.820
1124.000000000,-0.16243,-594.00,-1718.8,-84.017,-466.55,-9.0353,-18.708
1125.000000000,-0.16226,-593.11,-1717.8,-84.011,-466.36,-9.0297,-18.666
1126.000000000,-0.16215,-592.34,-1717.0,-84.005,-466.21,-9.0257,-18.640
1127.000000000,-0.16208,-591.65,-1716.2,-84.000,-466.10,-9.0229,-18.622
1128.000000000,-0.16203,-591.01,-1715.5,-83.994,-466.01,-9.0210,-18.609
1129.000000000,-0.16200,-590.41,-1714.8,-83.989,-465.94,-9.0197,-18.599
1130.000000000,-0.16198,-589.85,-1714.1,-83.983,-465.89,-9.0188,-18.592
1131.000000000,-0.16196,-589.31,-1713.4,-83.977,-465.84,-9.0180,-18.586
1132.000000000,-0.16194,-588.79,-1712.8,-83.971,-465.81,-9.0175,-18.582
1133.000000000,-0.16193,-588.29,-1712.2,-83.966,-465.78,-9.0171,-18.579
1134.000000000,-0.16192,-587.80,-1711.6,-83.960,-465.75,-9.0167,-18.576
1135.000000000,-0.16190,-587.30,-1711.0,-83.955,-465.72,-9.0164,-18.574
1136.000000000,-0.16189,-586.82,-1710.4,-83.950,-465.70,-9.0161,-18.572
1137.000000000,-0.16189,-586.34,-1709.8,-83.946,-465.68,-9.0158,-18.570
1138.000000000,-0.16188,-585.87,-1709.3,-83.941,-465.67,-9.0156,-18.569
1139.000000000,-0.16187,-585.42,-1708.7,-83.936,-465.65,-9.0154,-18.568
1140.000000000,-0.16186,-584.97,-1708.2,-83.931,-465.63,-9.0151,-18.567
1141.000000000,-0.16185,-584.54,-1707.7,-83.927,-465.62,-9.0149,-18.566
1142.000000000,-0.16184,-584.12,-1707.1,-83.922,-465.60,-9.0146,-18.565
1143.000000000,-0.16183,-583.71,-1706.6,-83.917,-465.59,-9.0144,-18.565
1144.000000000,-0.16182,-583.30,-1706.1,-83.913,-465.58,-9.0142,-18.564
1145.000000000,-0.16182,-582.90,-1705.5,-83.908,-465.56,-9.0140,-18.563
1146.000000000,-0.16181,-582.52,-1705.0,-83.904,-465.55,-9.0137,-18.563
1147.000000000,-0.16180,-582.12,-1704.5,-83.899,-465.54,-9.0135,-18.562
1148.000000000,-0.16214,1977.4,4078.5,-53.961,-371.64,-9.0262,-19.156
1149.000000000,-0.16301,1973.5,4074.4,-53.967,-372.83,-9.0565,-20.299
1150.000000000,-0.16270,-588.84,-1711.7,-83.904,-467.09,-9.0458,-18.877
1151.000000000,-0.16236,-587.43,-1710.1,-83.896,-466.53,-9.0360,-18.743
1152.000000000,-0.16214,-586.38,-1708.9,-83.892,-466.28,-9.0285,-18.689
1153.000000000,-0.16200,-585.52,-1707.9,-83.888,-466.08,-9.0233,-18.655
1154.000000000,-0.16192,-584.77,-1707.0,-83.884,-465.93,-9.0197,-18.631
1155.000000000,-0.16187,-584.15,-1706.2,-83.880,-465.82,-9.0173,-18.614
1156.000000000,-0.16183,-583.59,-1705.4,-83.877,-465.73,-9.0156,-18.601
1157.000000000,-0.16181,-583.03,-1704.7,-83.873,-465.66,-9.0143,-18.591
1158.000000000,-0.16179,-582.51,-1704.0,-83.869,-465.60,-9.0134,-18.584
1159.000000000,-0.16177,-582.03,-1703.3,-83.865,-465.56,-9.0128,-18.578
1160.000000000,-0.16177,-581.55,-1702.6,-83.862,-465.52,-9.0122,-18.574
1161.000000000,-0.16176,-581.09,-1702.0,-83.858,-465.49,-9.0118,-18.570
1162.000000000,-0.16175,-580.65,-1701.4,-83.854,-465.46,-9.0114,-18.567
1163.000000000,-0.16334,1978.9,4081.7,-53.916,-372.56,-9.0668,-21.303
1164.000000000,-0.16399,1975.1,4077.7,-53.923,-373.90,-9.0897,-20.739
1165.000000000,-0.16483,1971.9,4074.2,-53.926,-375.04,-9.1216,-21.675
1166.000000000,-0.16542,1968.6,4071.0,-53.930,-376.00,-9.1443,-21.869
1167.000000000,-0.16522,1964.4,4068.0,-53.937,-376.31,-9.1403,-21.004
1168.000000000,-0.16411,-595.91,-1717.2,-83.878,-469.82,-9.1033,-19.369
1169.000000000,-0.16328,-594.22,-1715.1,-83.875,-468.63,-9.0748,-19.103
1170.000000000,-0.16275,-592.95,-1713.5,-83.876,-467.89,-9.0548,-18.959
1171.000000000,-0.16243,-591.86,-1712.1,-83.878,-467.34,-9.0413,-18.861
1172.000000000,-0.16225,1968.2,4071.6,-53.944,-372.78,-9.0342,-18.839
1173.000000000,-0.16211,-594.28,-1714.3,-83.888,-467.03,-9.0271,-18.747
1174.000000000,-0.16276,1966.3,4069.9,-53.948,-372.88,-9.0489,-19.971
1175.000000000,-0.16253,-595.89,-1715.8,-83.890,-467.29,-9.0397,-18.876
1176.000000000,-0.16228,-594.23,-1713.9,-83.883,-466.70,-9.0317,-18.762
1177.000000000,-0.16211,-592.92,-1712.3,-83.880,-466.42,-9.0256,-18.710
1178.000000000,-0.16201,-591.80,-1711.0,-83.878,-466.21,-9.0214,-18.676
1179.000000000,-0.16204,1968.2,4072.7,-53.941,-371.97,-9.0228,-18.819
1180.000000000,-0.16198,-594.32,-1713.4,-83.883,-466.42,-9.0193,-18.660
1181.000000000,-0.16192,-593.00,-1711.8,-83.877,-465.98,-9.0171,-18.634
1182.000000000,-0.16188,-591.96,-1710.5,-83.873,-465.86,-9.0154,-18.618
1183.000000000,-0.16185,-591.04,-1709.3,-83.870,-465.77,-9.0141,-18.607
1184.000000000,-0.16183,-590.24,-1708.2,-83.865,-465.70,-9.0132,-18.598
1185.000000000,-0.16182,-589.54,-1707.2,-83.861,-465.65,-9.0125,-18.592
1186.000000000,-0.16181,-588.89,-1706.3,-83.855,-465.61,-9.0120,-18.587
1187.000000000,-0.16182,1970.8,4077.1,-53.916,-371.42,-9.0132,-18.611
1188.000000000,-0.16181,-591.95,-1709.3,-83.857,-465.95,-9.0120,-18.585
1189.000000000,-0.16180,-590.75,-1707.9,-83.849,-465.60,-9.0115,-18.580
1190.000000000,-0.16179,-589.81,-1706.7,-83.843,-465.55,-9.0111,-18.577
1191.000000000,-0.16178,-589.03,-1705.7,-83.838,-465.51,-9.0108,-18.575
1192.000000000,-0.16177,-588.30,-1704.8,-83.833,-465.49,-9.0105,-18.573
1193.000000000,-0.16176,-587.62,-1703.9,-83.828,-465.46,-9.0102,-18.571
1194.000000000,-0.16175,-586.98,-1703.1,-83.823,-465.44,-9.0100,-18.570
1195.000000000,-0.16175,-586.38,-1702.3,-83.818,-465.42,-9.0098,-18.569
1196.000000000,-0.16174,-585.81,-1701.6,-83.814,-465.41,-9.0096,-18.568
1197.000000000,-0.16176,1973.9,4081.6,-53.874,-371.26,-9.0113,-18.612
1198.000000000,-0.16175,-588.95,-1704.9,-83.815,-465.80,-9.0101,-18.574
1199.000000000,-0.16240,1971.3,4078.9,-53.872,-371.83,-9.0333,-19.703
1200.000000000,-0.16224,-591.11,-1707.2,-83.811,-466.40,-9.0274,-18.750
1201.000000000,-0.16205,-589.70,-1705.6,-83.803,-465.96,-9.0219,-18.668
1202.000000000,-0.16192,-588.59,-1704.4,-83.797,-465.80,-9.0176,-18.636
1203.000000000,-0.16621,1971.5,4079.2,-53.859,-375.02,-9.1652,-26.121
1204.000000000,-0.16614,1967.5,4075.3,-53.867,-376.52,-9.1642,-21.451
1205.000000000,-0.16471,1962.8,4072.1,-53.874,-376.02,-9.1230,-19.562
1206.000000000,-0.16365,1959.6,4069.1,-53.881,-375.19,-9.0893,-19.243
1207.000000000,-0.16298,-600.00,-1716.0,-83.822,-468.61,-9.0636,-19.043
1208.000000000,-0.16256,-598.20,-1713.9,-83.820,-467.63,-9.0469,-18.941
1209.000000000,-0.16229,-596.75,-1712.2,-83.821,-467.11,-9.0353,-18.834
1210.000000000,-0.16219,1963.5,4071.8,-53.886,-372.62,-9.0309,-18.890
1211.000000000,-0.16206,-598.71,-1713.9,-83.830,-466.90,-9.0243,-18.745
1212.000000000,-0.16197,-597.10,-1712.0,-83.825,-466.34,-9.0200,-18.701
1213.000000000,-0.16234,1963.3,4072.1,-53.888,-372.32,-9.0329,-19.416
1214.000000000,-0.16220,-598.91,-1713.7,-83.830,-466.76,-9.0268,-18.769
1215.000000000,-0.16205,-597.28,-1711.8,-83.824,-466.26,-9.0218,-18.699
1216.000000000,-0.16197,-595.97,-1710.2,-83.822,-466.07,-9.0185,-18.688
1217.000000000,-0.16190,-594.89,-1708.9,-83.820,-465.93,-9.0157,-18.647
1218.000000000,-0.16187,1965.2,4074.8,-53.883,-371.67,-9.0154,-18.658
1219.000000000,-0.16184,-597.34,-1711.2,-83.825,-466.15,-9.0131,-18.621
1220.000000000,-0.16182,-595.94,-1709.5,-83.818,-465.74,-9.0119,-18.609
1221.000000000,-0.16180,-594.81,-1708.1,-83.814,-465.66,-9.0110,-18.601
1222.000000000,-0.16179,-593.85,-1706.9,-83.810,-465.60,-9.0103,-18.595
1223.000000000,-0.16178,-593.01,-1705.8,-83.806,-465.55,-9.0098,-18.590
1224.000000000,-0.16177,-592.24,-1704.8,-83.801,-465.52,-9.0094,-18.586
1225.000000000,-0.16191,1967.6,4078.7,-53.863,-371.44,-9.0150,-18.827
1226.000000000,-0.16187,-595.03,-1707.6,-83.805,-465.99,-9.0130,-18.620
1227.000000000,-0.16183,-593.70,-1706.1,-83.797,-465.62,-9.0116,-18.600
1228.000000000,-0.16180,-592.64,-1704.9,-83.792,-465.55,-9.0105,-18.592
1229.000000000,-0.16180,1967.4,4078.6,-53.854,-371.35,-9.0113,-18.618
1230.000000000,-0.16178,-595.16,-1707.5,-83.794,-465.88,-9.0099,-18.591
1231.000000000,-0.16199,1965.3,4076.5,-53.852,-371.54,-9.0180,-18.973
1232.000000000,-0.16207,1961.3,4073.1,-53.859,-372.02,-9.0210,-18.887
1233.000000000,-0.16197,-599.38,-1712.3,-83.796,-466.19,-9.0171,-18.659
1234.000000000,-0.16241,1961.1,4072.2,-53.854,-372.02,-9.0334,-19.533
1235.000000000,-0.16362,1957.1,4069.2,-53.859,-373.46,-9.0750,-21.132
1236.000000000,-0.16340,1954.8,4066.7,-53.862,-373.73,-9.0689,-19.535
1237.000000000,-0.16284,-604.37,-1718.2,-83.800,-467.61,-9.0510,-18.934
1238.000000000,-0.16243,-602.33,-1715.8,-83.793,-466.86,-9.0374,-18.816
1239.000000000,-0.16218,-600.64,-1713.9,-83.790,-466.49,-9.0279,-18.750
1240.000000000,-0.16203,-599.21,-1712.2,-83.787,-466.21,-9.0213,-18.704
1241.000000000,-0.16193,-597.94,-1710.7,-83.784,-466.01,-9.0170,-18.672
1242.000000000,-0.16186,-596.78,-1709.3,-83.781,-465.85,-9.0139,-18.648
1243.000000000,-0.16183,-595.72,-1708.1,-83.778,-465.74,-9.0123,-18.651
1244.000000000,-0.16180,-594.74,-1707.0,-83.775,-465.64,-9.0107,-18.620
1245.000000000,-0.16178,-593.83,-1705.9,-83.773,-465.57,-9.0095,-18.608
1246.000000000,-0.16183,1966.1,4077.5,-53.835,-371.40,-9.0118,-18.707
1247.000000000,-0.16180,-596.40,-1708.7,-83.777,-465.92,-9.0100,-18.611
1248.000000000,-0.16193,1964.1,4075.4,-53.836,-371.51,-9.0154,-18.870
1249.000000000,-0.16472,1959.9,4072.0,-53.843,-374.12,-9.1109,-23.510
1250.000000000,-0.16465,1956.6,4069.1,-53.846,-374.90,-9.1098,-20.459
1251.000000000,-0.16375,1953.8,4066.4,-53.851,-374.58,-9.0841,-19.300
1252.000000000,-0.16303,-605.27,-1718.5,-83.789,-468.18,-9.0600,-19.003
1253.000000000,-0.16257,-603.24,-1716.1,-83.783,-467.27,-9.0431,-18.882
1254.000000000,-0.16229,-601.60,-1714.1,-83.780,-466.80,-9.0316,-18.802
1255.000000000,-0.16211,-600.24,-1712.5,-83.779,-466.46,-9.0239,-18.746
1256.000000000,-0.16200,-599.03,-1711.1,-83.779,-466.21,-9.0188,-18.706
1257.000000000,-0.16192,-597.90,-1709.7,-83.777,-466.01,-9.0152,-18.675
1258.000000000,-0.16187,-596.86,-1708.4,-83.774,-465.86,-9.0128,-18.652
1259.000000000,-0.16184,-595.85,-1707.2,-83.771,-465.74,-9.0111,-18.635
1260.000000000,-0.16184,1964.2,4076.4,-53.833,-371.52,-9.0120,-18.673
1261.000000000,-0.16182,-598.21,-1709.7,-83.774,-466.01,-9.0101,-18.620
1262.000000000,-0.16179,-596.71,-1708.0,-83.766,-465.62,-9.0092,-18.608
1263.000000000,-0.16178,-595.46,-1706.7,-83.762,-465.53,-9.0084,-18.600
1264.000000000,-0.16176,-594.39,-1705.5,-83.758,-465.48,-9.0078,-18.594
1265.000000000,-0.16175,-593.44,-1704.4,-83.754,-465.43,-9.0074,-18.589
1266.000000000,-0.16174,-592.59,-1703.4,-83.749,-465.40,-9.0070,-18.586
1267.000000000,-0.16236,1967.3,4080.1,-53.810,-371.72,-9.0293,-19.662
1268.000000000,-0.16222,-595.31,-1706.1,-83.751,-466.31,-9.0237,-18.754
1269.000000000,-0.16204,-593.99,-1704.7,-83.743,-465.87,-9.0186,-18.674
1270.000000000,-0.16192,-592.91,-1703.4,-83.738,-465.72,-9.0145,-18.644
1271.000000000,-0.16184,-591.97,-1702.3,-83.733,-465.61,-9.0117,-18.625
1272.000000000,-0.16179,-591.11,-1701.3,-83.729,-465.52,-9.0097,-18.611
1273.000000000,-0.16237,1968.8,4082.1,-53.790,-371.78,-9.0302,-19.643
1274.000000000,-0.16696,1965.3,4078.4,-53.796,-375.99,-9.1876,-26.914
1275.000000000,-0.16588,1959.8,4074.7,-53.804,-376.53,-9.1532,-20.271
1276.000000000,-0.16446,1956.4,4071.8,-53.811,-375.84,-9.1132,-19.507
1277.000000000,-0.16347,-602.90,-1713.4,-83.752,-469.14,-9.0794,-19.172
1278.000000000,-0.16285,-601.09,-1711.4,-83.750,-468.02,-9.0562,-19.016
1279.000000000,-0.16246,-599.55,-1709.6,-83.749,-467.39,-9.0406,-18.901
1280.000000000,-0.16222,-598.24,-1708.0,-83.748,-466.92,-9.0301,-18.823
1281.000000000,-0.16206,-597.10,-1706.6,-83.747,-466.57,-9.0231,-18.766
1282.000000000,-0.16195,-596.08,-1705.3,-83.746,-466.30,-9.0183,-18.723
1283.000000000,-0.16188,-595.11,-1704.1,-83.743,-466.10,-9.0150,-18.691
1284.000000000,-0.16183,-594.21,-1703.0,-83.741,-465.94,-9.0127,-18.666
1285.000000000,-0.16179,-593.37,-1701.9,-83.740,-465.82,-9.0110,-18.647
1286.000000000,-0.16176,-592.64,-1701.0,-83.738,-465.72,-9.0098,-18.633
1287.000000000,-0.16175,-591.98,-1700.1,-83.736,-465.65,-9.0091,-18.631
1288.000000000,-0.16173,-591.36,-1699.2,-83.735,-465.58,-9.0084,-18.614
1289.000000000,-0.16172,-590.80,-1698.4,-83.732,-465.53,-9.0078,-18.606
1290.000000000,-0.16170,-590.29,-1697.6,-83.729,-465.49,-9.0073,-18.601
1291.000000000,-0.16169,-589.77,-1696.8,-83.726,-465.46,-9.0070,-18.596
1292.000000000,-0.16168,-589.20,-1696.1,-83.723,-465.43,-9.0067,-18.592
1293.000000000,-0.16168,-588.65,-1695.4,-83.720,-465.40,-9.0064,-18.590
1294.000000000,-0.16167,-588.12,-1694.7,-83.717,-465.38,-9.0062,-18.587
1295.000000000,-0.16166,-587.57,-1694.1,-83.715,-465.36,-9.0060,-18.585
1296.000000000,-0.16166,-587.02,-1693.5,-83.713,-465.35,-9.0058,-18.584
1297.000000000,-0.16165,-586.48,-1692.8,-83.711,-465.33,-9.0057,-18.582
1298.000000000,-0.16164,-585.96,-1692.2,-83.709,-465.32,-9.0055,-18.581
1299.000000000,-0.16164,-585.44,-1691.6,-83.707,-465.30,-9.0053,-18.580
1300.000000000,-0.16163,-584.97,-1691.0,-83.705,-465.29,-9.0052,-18.579
1301.000000000,-0.16163,-584.52,-1690.4,-83.702,-465.28,-9.0050,-18.578
1302.000000000,-0.16162,-584.07,-1689.9,-83.700,-465.27,-9.0049,-18.578
1303.000000000,-0.16164,1975.5,4093.2,-53.764,-371.11,-9.0064,-18.605
1304.000000000,-0.16214,1971.7,4089.1,-53.773,-371.90,-9.0234,-19.432
1305.000000000,-0.16207,1968.2,4085.6,-53.779,-372.04,-9.0213,-18.795
1306.000000000,-0.16192,-593.29,-1699.9,-83.717,-466.16,-9.0162,-18.667
1307.000000000,-0.16184,1967.4,4084.4,-53.774,-371.55,-9.0143,-18.673
1308.000000000,-0.16176,-594.34,-1701.2,-83.715,-465.97,-9.0108,-18.626
1309.000000000,-0.16171,-592.56,-1699.4,-83.707,-465.55,-9.0087,-18.612
1310.000000000,-0.16167,-591.14,-1697.9,-83.702,-465.44,-9.0073,-18.602
1311.000000000,-0.16165,-589.95,-1696.6,-83.698,-465.37,-9.0063,-18.595
1312.000000000,-0.16163,-588.91,-1695.5,-83.693,-465.32,-9.0055,-18.589
1313.000000000,-0.16161,-588.00,-1694.5,-83.689,-465.28,-9.0049,-18.585
1314.000000000,-0.16160,-587.20,-1693.6,-83.685,-465.25,-9.0045,-18.582
1315.000000000,-0.16159,-586.45,-1692.7,-83.681,-465.22,-9.0041,-18.579
1316.000000000,-0.16158,-585.78,-1691.9,-83.676,-465.19,-9.0038,-18.577
1317.000000000,-0.16157,-585.16,-1691.1,-83.671,-465.17,-9.0036,-18.576
1318.000000000,-0.16156,-584.56,-1690.4,-83.667,-465.15,-9.0033,-18.574
1319.000000000,-0.16156,-583.97,-1689.7,-83.662,-465.14,-9.0031,-18.573
1320.000000000,-0.16155,-583.39,-1689.0,-83.658,-465.12,-9.0029,-18.572
1321.000000000,-0.16328,1976.3,4094.2,-53.719,-372.34,-9.0635,-21.563
1322.000000000,-0.16440,1972.6,4090.2,-53.725,-374.10,-9.1024,-21.636
1323.000000000,-0.16415,1969.6,4086.9,-53.727,-374.52,-9.0976,-20.236
1324.000000000,-0.16340,1965.6,4083.8,-53.732,-374.21,-9.0753,-19.340
1325.000000000,-0.16381,1962.7,4081.0,-53.737,-374.53,-9.0901,-20.807
1326.000000000,-0.16347,1960.3,4078.5,-53.741,-374.41,-9.0781,-19.721
1327.000000000,-0.16297,1958.0,4076.1,-53.746,-374.01,-9.0612,-19.261
1328.000000000,-0.16615,1955.9,4073.8,-53.752,-376.45,-9.1697,-25.223
1329.000000000,-0.16548,1952.9,4071.3,-53.763,-376.75,-9.1465,-20.631
1330.000000000,-0.16488,1950.3,4068.8,-53.777,-376.53,-9.1307,-20.669
1331.000000000,-0.16467,1948.2,4066.6,-53.792,-376.40,-9.1243,-20.866
1332.000000000,-0.16371,-609.93,-1717.8,-83.736,-469.79,-9.0898,-19.369
1333.000000000,-0.16310,1948.9,4067.6,-53.801,-374.51,-9.0689,-19.319
1334.000000000,-0.16262,-609.91,-1717.1,-83.745,-468.33,-9.0492,-19.015
1335.000000000,-0.16229,-607.84,-1714.4,-83.743,-467.43,-9.0359,-18.905
1336.000000000,-0.16215,1951.1,4070.3,-53.810,-372.85,-9.0300,-18.932
1337.000000000,-0.16226,1947.6,4067.6,-53.821,-373.11,-9.0328,-19.246
1338.000000000,-0.16222,1945.1,4065.3,-53.828,-373.03,-9.0304,-19.018
1339.000000000,-0.16230,1943.0,4063.4,-53.832,-373.03,-9.0329,-19.209
1340.000000000,-0.16226,1941.1,4061.5,-53.836,-372.98,-9.0314,-19.050
1341.000000000,-0.16222,1939.3,4059.8,-53.840,-372.91,-9.0301,-19.028
1342.000000000,-0.16257,1937.5,4058.2,-53.843,-373.16,-9.0421,-19.668
1343.000000000,-0.16233,-619.79,-1726.0,-83.781,-467.20,-9.0328,-18.872
1344.000000000,-0.16210,-617.15,-1722.9,-83.773,-466.58,-9.0251,-18.765
1345.000000000,-0.16195,-615.29,-1720.3,-83.769,-466.31,-9.0194,-18.726
1346.000000000,-0.16185,-613.70,-1718.2,-83.767,-466.11,-9.0154,-18.688
1347.000000000,-0.16178,-612.22,-1716.3,-83.764,-465.96,-9.0125,-18.665
1348.000000000,-0.16174,-610.89,-1714.6,-83.761,-465.84,-9.0106,-18.649
1349.000000000,-0.16171,-609.61,-1713.0,-83.758,-465.75,-9.0092,-18.636
1350.000000000,-0.16188,1948.6,4071.0,-53.821,-371.66,-9.0156,-18.945
1351.000000000,-0.16182,-611.33,-1714.8,-83.762,-466.18,-9.0127,-18.670
1352.000000000,-0.16224,1946.6,4069.5,-53.821,-372.01,-9.0281,-19.465
1353.000000000,-0.16214,1943.5,4066.4,-53.829,-372.40,-9.0248,-18.838
1354.000000000,-0.16218,1941.2,4063.8,-53.835,-372.51,-9.0272,-19.072
1355.000000000,-0.16202,-616.53,-1721.1,-83.774,-466.59,-9.0207,-18.731
1356.000000000,-0.16189,-614.27,-1718.6,-83.768,-466.08,-9.0160,-18.684
1357.000000000,-0.16181,-612.52,-1716.5,-83.765,-465.90,-9.0127,-18.659
1358.000000000,-0.16175,-611.00,-1714.7,-83.763,-465.78,-9.0103,-18.642
1359.000000000,-0.16172,-609.65,-1713.1,-83.761,-465.69,-9.0086,-18.630
1360.000000000,-0.16170,-608.43,-1711.7,-83.758,-465.61,-9.0075,-18.621
1361.000000000,-0.16169,-607.29,-1710.3,-83.755,-465.56,-9.0067,-18.614
1362.000000000,-0.16168,-606.21,-1709.1,-83.752,-465.51,-9.0061,-18.608
1363.000000000,-0.16168,-605.18,-1707.9,-83.749,-465.48,-9.0057,-18.604
1364.000000000,-0.16397,1953.5,4075.7,-53.810,-373.13,-9.0851,-22.548
1365.000000000,-0.16873,1948.7,4072.0,-53.817,-377.96,-9.2490,-28.297
1366.000000000,-0.16749,1943.9,4068.2,-53.832,-378.68,-9.2124,-21.385
1367.000000000,-0.16549,-614.87,-1717.5,-83.782,-471.83,-9.1526,-19.796
1368.000000000,-0.16412,-613.14,-1715.7,-83.786,-470.22,-9.1069,-19.417
1369.000000000,-0.16327,-611.74,-1714.0,-83.789,-469.14,-9.0751,-19.197
1370.000000000,-0.16275,-610.55,-1712.4,-83.789,-468.31,-9.0537,-19.046
1371.000000000,-0.16242,-609.45,-1711.0,-83.788,-467.69,-9.0394,-18.939
1372.000000000,-0.16221,-608.41,-1709.7,-83.790,-467.22,-9.0298,-18.860
1373.000000000,-0.16207,-607.65,-1708.6,-83.790,-466.87,-9.0234,-18.801
1374.000000000,-0.16198,-607.00,-1707.5,-83.789,-466.60,-9.0191,-18.757
1375.000000000,-0.16192,-606.34,-1706.4,-83.787,-466.39,-9.0160,-18.723
1376.000000000,-0.16188,-605.73,-1705.4,-83.784,-466.22,-9.0138,-18.697
1377.000000000,-0.16186,-605.11,-1704.5,-83.781,-466.10,-9.0126,-18.697
1378.000000000,-0.16183,-604.51,-1703.6,-83.779,-466.00,-9.0114,-18.664
1379.000000000,-0.16181,-603.90,-1702.7,-83.776,-465.92,-9.0105,-18.651
1380.000000000,-0.16180,-603.33,-1701.9,-83.773,-465.85,-9.0098,-18.641
1381.000000000,-0.16178,-602.74,-1701.1,-83.770,-465.80,-9.0092,-18.633
1382.000000000,-0.16178,-602.12,-1700.3,-83.768,-465.75,-9.0088,-18.627
1383.000000000,-0.16177,-601.49,-1699.6,-83.766,-465.72,-9.0085,-18.622
1384.000000000,-0.16176,-600.87,-1698.9,-83.765,-465.68,-9.0082,-18.618
1385.000000000,-0.16176,-600.27,-1698.2,-83.763,-465.66,-9.0079,-18.615
1386.000000000,-0.16175,-599.70,-1697.6,-83.762,-465.64,-9.0077,-18.613
1387.000000000,-0.16175,-599.14,-1697.0,-83.762,-465.62,-9.0075,-18.611
1388.000000000,-0.16175,-598.62,-1696.4,-83.762,-465.60,-9.0074,-18.609
1389.000000000,-0.16175,-598.09,-1695.8,-83.761,-465.58,-9.0072,-18.607
1390.000000000,-0.16176,-597.55,-1695.2,-83.760,-465.58,-9.0074,-18.623
1391.000000000,-0.16176,-597.00,-1694.6,-83.759,-465.56,-9.0072,-18.608
1392.000000000,-0.16176,-596.45,-1694.0,-83.757,-465.55,-9.0070,-18.605
1393.000000000,-0.16176,-595.90,-1693.5,-83.754,-465.53,-9.0069,-18.604
1394.000000000,-0.16176,-595.35,-1692.9,-83.752,-465.52,-9.0067,-18.603
1395.000000000,-0.16176,-594.78,-1692.4,-83.749,-465.51,-9.0066,-18.602
1396.000000000,-0.16176,-594.22,-1691.9,-83.747,-465.50,-9.0065,-18.601
1397.000000000,-0.16175,-593.67,-1691.3,-83.745,-465.49,-9.0064,-18.601
1398.000000000,-0.16175,-593.13,-1690.8,-83.741,-465.47,-9.0062,-18.600
1399.000000000,-0.16175,-592.60,-1690.3,-83.737,-465.46,-9.0061,-18.599
1400.000000000,-0.16175,-592.06,-1689.8,-83.733,-465.45,-9.0060,-18.599
1401.000000000,-0.16174,-591.54,-1689.3,-83.730,-465.44,-9.0059,-18.598
1402.000000000,-0.16174,-591.04,-1688.8,-83.726,-465.43,-9.0058,-18.597
1403.000000000,-0.16174,-590.57,-1688.4,-83.722,-465.42,-9.0056,-18.597
1404.000000000,-0.16274,1969.0,4094.6,-53.784,-372.06,-9.0411,-20.329
1405.000000000,-0.16256,1965.0,4090.4,-53.791,-372.57,-9.0351,-18.936
1406.000000000,-0.16229,1960.3,4086.9,-53.794,-372.51,-9.0278,-18.790
1407.000000000,-0.16223,1957.5,4083.7,-53.797,-372.48,-9.0260,-18.947
1408.000000000,-0.16207,-601.85,-1701.6,-83.733,-466.52,-9.0195,-18.719
1409.000000000,-0.16195,-599.91,-1699.6,-83.726,-466.00,-9.0150,-18.680
1410.000000000,-0.16339,1960.4,4084.5,-53.787,-372.88,-9.0648,-21.259
1411.000000000,-0.16305,1955.8,4081.2,-53.794,-373.35,-9.0534,-19.139
1412.000000000,-0.16259,-603.57,-1704.2,-83.731,-467.28,-9.0390,-18.874
1413.000000000,-0.16228,-601.73,-1702.2,-83.724,-466.60,-9.0284,-18.790
1414.000000000,-0.16209,-600.21,-1700.6,-83.721,-466.29,-9.0209,-18.739
1415.000000000,-0.16196,-598.86,-1699.3,-83.717,-466.06,-9.0158,-18.703
1416.000000000,-0.16188,-597.67,-1698.1,-83.713,-465.89,-9.0124,-18.677
1417.000000000,-0.16183,-596.61,-1697.0,-83.709,-465.76,-9.0100,-18.658
1418.000000000,-0.16179,-595.62,-1696.0,-83.705,-465.66,-9.0083,-18.643
1419.000000000,-0.16177,-594.69,-1695.0,-83.701,-465.58,-9.0071,-18.632
1420.000000000,-0.16175,-593.79,-1694.1,-83.697,-465.51,-9.0062,-18.624
1421.000000000,-0.16173,-592.94,-1693.3,-83.692,-465.46,-9.0056,-18.617
1422.000000000,-0.16173,-592.14,-1692.4,-83.688,-465.42,-9.0050,-18.612
1423.000000000,-0.16172,-591.37,-1691.7,-83.683,-465.38,-9.0046,-18.608
1424.000000000,-0.16172,-590.62,-1690.9,-83.679,-465.36,-9.0043,-18.604
1425.000000000,-0.16171,-589.93,-1690.2,-83.675,-465.33,-9.0039,-18.602
1426.000000000,-0.16184,1969.8,4092.9,-53.736,-371.26,-9.0094,-18.836
1427.000000000,-0.16181,-592.86,-1693.5,-83.676,-465.81,-9.0075,-18.636
1428.000000000,-0.16176,-591.58,-1692.3,-83.668,-465.45,-9.0061,-18.618
1429.000000000,-0.16173,-590.53,-1691.3,-83.664,-465.38,-9.0050,-18.610
1430.000000000,-0.16171,-589.61,-1690.3,-83.659,-465.33,-9.0042,-18.605
1431.000000000,-0.16170,-588.76,-1689.5,-83.654,-465.30,-9.0036,-18.601
1432.000000000,-0.16169,-587.97,-1688.7,-83.649,-465.27,-9.0031,-18.598
1433.000000000,-0.16226,1971.9,4094.5,-53.710,-371.55,-9.0236,-19.592
1434.000000000,-0.16310,1968.4,4090.6,-53.716,-372.77,-9.0529,-20.440
1435.000000000,-0.16601,1965.5,4087.2,-53.719,-375.47,-9.1541,-24.614
1436.000000000,-0.16522,1961.6,4084.0,-53.723,-375.85,-9.1298,-20.263
1437.000000000,-0.16399,-599.30,-1701.4,-83.662,-469.36,-9.0926,-19.329
1438.000000000,-0.16315,-597.35,-1699.3,-83.656,-468.20,-9.0643,-19.099
1439.000000000,-0.16263,-595.85,-1697.7,-83.654,-467.51,-9.0446,-18.963
1440.000000000,-0.16231,-594.63,-1696.4,-83.653,-466.98,-9.0313,-18.870
1441.000000000,-0.16211,-593.55,-1695.2,-83.652,-466.59,-9.0224,-18.804
1442.000000000,-0.16198,-592.55,-1694.1,-83.649,-466.29,-9.0164,-18.755
1443.000000000,-0.16197,1967.5,4089.5,-53.712,-371.96,-9.0161,-18.855
1444.000000000,-0.16190,-595.00,-1696.7,-83.654,-466.35,-9.0119,-18.713
1445.000000000,-0.16184,-593.57,-1695.1,-83.647,-465.88,-9.0093,-18.682
1446.000000000,-0.16182,-592.40,-1693.8,-83.642,-465.74,-9.0078,-18.688
1447.000000000,-0.16179,-591.41,-1692.7,-83.638,-465.64,-9.0063,-18.651
1448.000000000,-0.16177,-590.51,-1691.6,-83.633,-465.55,-9.0052,-18.638
1449.000000000,-0.16175,-589.68,-1690.6,-83.629,-465.48,-9.0043,-18.629
1450.000000000,-0.16174,-588.91,-1689.8,-83.624,-465.43,-9.0036,-18.621
1451.000000000,-0.16173,-588.19,-1689.0,-83.620,-465.39,-9.0031,-18.616
1452.000000000,-0.16180,1971.6,4094.5,-53.681,-371.25,-9.0063,-18.743
1453.000000000,-0.16177,-591.11,-1691.9,-83.621,-465.79,-9.0047,-18.629
1454.000000000,-0.16188,1969.2,4091.9,-53.678,-371.37,-9.0094,-18.850
1455.000000000,-0.16183,-593.11,-1694.1,-83.617,-465.88,-9.0069,-18.649
1456.000000000,-0.16178,-591.62,-1692.5,-83.608,-465.49,-9.0052,-18.628
1457.000000000,-0.16174,-590.45,-1691.3,-83.602,-465.41,-9.0039,-18.618
1458.000000000,-0.16172,-589.45,-1690.3,-83.596,-465.35,-9.0029,-18.612
1459.000000000,-0.16170,-588.56,-1689.3,-83.591,-465.31,-9.0022,-18.607
1460.000000000,-0.16172,1971.4,4094.6,-53.651,-371.14,-9.0038,-18.662
1461.000000000,-0.16171,-591.22,-1692.1,-83.591,-465.68,-9.0026,-18.620
1462.000000000,-0.16169,-589.87,-1690.7,-83.582,-465.33,-9.0019,-18.607
1463.000000000,-0.16176,1970.3,4093.4,-53.641,-371.18,-9.0052,-18.742
1464.000000000,-0.16173,-592.09,-1693.1,-83.581,-465.71,-9.0034,-18.622
1465.000000000,-0.16170,-590.60,-1691.7,-83.572,-465.34,-9.0023,-18.610
1466.000000000,-0.16167,-589.41,-1690.5,-83.566,-465.28,-9.0014,-18.604
1467.000000000,-0.16166,-588.35,-1689.4,-83.562,-465.23,-9.0008,-18.600
1468.000000000,-0.16165,-587.41,-1688.5,-83.557,-465.20,-9.0002,-18.598
1469.000000000,-0.16164,-586.55,-1687.7,-83.552,-465.18,-8.9998,-18.595
1470.000000000,-0.16163,-585.75,-1686.9,-83.547,-465.16,-8.9995,-18.594
1471.000000000,-0.16162,-585.00,-1686.1,-83.542,-465.14,-8.9992,-18.592
1472.000000000,-0.16161,-584.29,-1685.4,-83.537,-465.12,-8.9990,-18.591
1473.000000000,-0.16161,-583.62,-1684.7,-83.532,-465.11,-8.9987,-18.590
1474.000000000,-0.16160,-582.97,-1684.1,-83.527,-465.09,-8.9985,-18.589
1475.000000000,-0.16172,1976.8,4099.8,-53.588,-371.02,-9.0036,-18.804
1476.000000000,-0.16194,1973.1,4096.1,-53.594,-371.62,-9.0113,-19.049
1477.000000000,-0.16239,1970.1,4092.9,-53.597,-372.12,-9.0272,-19.611
1478.000000000,-0.16218,-591.61,-1693.1,-83.534,-466.31,-9.0195,-18.789
1479.000000000,-0.16266,1969.4,4091.9,-53.591,-372.19,-9.0378,-19.899
1480.000000000,-0.16237,-592.49,-1694.2,-83.531,-466.62,-9.0270,-18.862
1481.000000000,-0.16210,-590.62,-1692.4,-83.524,-466.05,-9.0182,-18.754
1482.000000000,-0.16192,-589.14,-1690.9,-83.519,-465.80,-9.0116,-18.706
1483.000000000,-0.16180,-587.94,-1689.7,-83.514,-465.61,-9.0070,-18.675
1484.000000000,-0.16173,-586.89,-1688.5,-83.510,-465.47,-9.0039,-18.653
1485.000000000,-0.16169,-585.92,-1687.5,-83.506,-465.36,-9.0017,-18.636
1486.000000000,-0.16165,-585.03,-1686.6,-83.502,-465.28,-9.0002,-18.624
1487.000000000,-0.16163,-584.19,-1685.7,-83.498,-465.21,-8.9992,-18.615
1488.000000000,-0.16162,-583.38,-1684.9,-83.493,-465.15,-8.9984,-18.608
1489.000000000,-0.16165,1976.5,4099.1,-53.554,-370.98,-9.0002,-18.671
1490.000000000,-0.16163,-586.11,-1687.8,-83.494,-465.51,-8.9987,-18.610
1491.000000000,-0.16161,-584.76,-1686.5,-83.486,-465.14,-8.9979,-18.601
1492.000000000,-0.16159,-583.67,-1685.5,-83.481,-465.08,-8.9973,-18.596
1493.000000000,-0.16158,-582.71,-1684.6,-83.476,-465.04,-8.9969,-18.593
1494.000000000,-0.16157,-581.85,-1683.8,-83.471,-465.01,-8.9965,-18.590
1495.000000000,-0.16156,-581.06,-1683.0,-83.467,-464.99,-8.9962,-18.588
1496.000000000,-0.16155,-580.31,-1682.3,-83.462,-464.97,-8.9959,-18.587
1497.000000000,-0.16157,1979.5,4101.6,-53.523,-370.81,-8.9975,-18.623
1498.000000000,-0.16156,-583.15,-1685.3,-83.464,-465.35,-8.9963,-18.591
1499.000000000,-0.16154,-581.86,-1684.1,-83.455,-465.00,-8.9959,-18.587
1500.000000000,-0.16153,-580.81,-1683.1,-83.450,-464.96,-8.9956,-18.585
1501.000000000,-0.16152,-579.90,-1682.3,-83.446,-464.93,-8.9953,-18.583
1502.000000000,-0.16152,-579.08,-1681.5,-83.441,-464.90,-8.9950,-18.582
1503.000000000,-0.16151,-578.31,-1680.7,-83.436,-464.88,-8.9948,-18.581
1504.000000000,-0.16150,-577.58,-1680.0,-83.431,-464.87,-8.9945,-18.580
1505.000000000,-0.16150,-576.88,-1679.4,-83.426,-464.85,-8.9944,-18.580
1506.000000000,-0.16373,1982.9,4104.5,-53.486,-372.47,-9.0720,-22.428
1507.000000000,-0.16322,-579.79,-1682.5,-83.426,-467.24,-9.0546,-19.193
1508.000000000,-0.16260,-578.54,-1681.3,-83.417,-466.58,-9.0370,-18.917
1509.000000000,-0.16223,1981.5,4102.8,-53.477,-372.05,-9.0259,-18.886
1510.000000000,-0.16196,-581.14,-1684.0,-83.419,-466.29,-9.0153,-18.763
1511.000000000,-0.16179,-579.76,-1682.7,-83.410,-465.70,-9.0085,-18.714
1512.000000000,-0.16198,1980.4,4101.7,-53.470,-371.55,-9.0151,-19.190
1513.000000000,-0.16184,-582.00,-1685.0,-83.411,-465.97,-9.0090,-18.738
1514.000000000,-0.16171,-580.56,-1683.6,-83.402,-465.48,-9.0045,-18.683
1515.000000000,-0.16162,-579.41,-1682.4,-83.397,-465.30,-9.0012,-18.656
1516.000000000,-0.16156,-578.44,-1681.4,-83.393,-465.17,-8.9988,-18.637
1517.000000000,-0.16152,-577.56,-1680.5,-83.388,-465.08,-8.9971,-18.623
1518.000000000,-0.16150,-576.74,-1679.6,-83.384,-465.00,-8.9959,-18.612
1519.000000000,-0.16147,-575.99,-1678.8,-83.379,-464.94,-8.9950,-18.604
1520.000000000,-0.16146,-575.30,-1678.1,-83.375,-464.89,-8.9944,-18.598
1521.000000000,-0.16144,-574.66,-1677.4,-83.371,-464.85,-8.9938,-18.593
1522.000000000,-0.16143,-574.06,-1676.8,-83.366,-464.82,-8.9934,-18.589
1523.000000000,-0.16142,-573.47,-1676.2,-83.362,-464.79,-8.9931,-18.586
1524.000000000,-0.16141,-572.91,-1675.7,-83.358,-464.77,-8.9928,-18.584
1525.000000000,-0.16156,1986.7,4108.4,-53.419,-370.71,-8.9989,-18.845
1526.000000000,-0.16152,-576.08,-1678.7,-83.360,-465.26,-8.9967,-18.623
1527.000000000,-0.16147,-574.93,-1677.5,-83.352,-464.89,-8.9953,-18.603
1528.000000000,-0.16143,-574.00,-1676.6,-83.347,-464.82,-8.9941,-18.594
1529.000000000,-0.16141,-573.20,-1675.9,-83.343,-464.78,-8.9933,-18.589
1530.000000000,-0.16139,-572.48,-1675.2,-83.338,-464.74,-8.9926,-18.585
1531.000000000,-0.16142,1987.3,4109.1,-53.399,-370.58,-8.9945,-18.648
1532.000000000,-0.16140,-575.42,-1677.9,-83.340,-465.12,-8.9931,-18.593
1533.000000000,-0.16138,-574.20,-1676.7,-83.332,-464.76,-8.9925,-18.584
1534.000000000,-0.16137,-573.23,-1675.8,-83.326,-464.71,-8.9920,-18.585
1535.000000000,-0.16135,-572.39,-1675.0,-83.322,-464.67,-8.9915,-18.579
1536.000000000,-0.16134,-571.65,-1674.3,-83.318,-464.65,-8.9911,-18.577
1537.000000000,-0.16133,-570.97,-1673.7,-83.313,-464.62,-8.9908,-18.575
1538.000000000,-0.16132,-570.34,-1673.1,-83.309,-464.60,-8.9905,-18.574
1539.000000000,-0.16132,-569.76,-1672.5,-83.305,-464.58,-8.9903,-18.573
1540.000000000,-0.16131,-569.21,-1672.0,-83.301,-464.57,-8.9900,-18.572
1541.000000000,-0.16130,-568.69,-1671.5,-83.296,-464.55,-8.9898,-18.571
1542.000000000,-0.16130,-568.20,-1671.0,-83.292,-464.54,-8.9896,-18.570
1543.000000000,-0.16129,-567.73,-1670.5,-83.287,-464.52,-8.9894,-18.569
1544.000000000,-0.16131,1991.8,4114.7,-53.348,-370.37,-8.9912,-18.615
1545.000000000,-0.16130,-571.05,-1673.4,-83.289,-464.92,-8.9901,-18.576
1546.000000000,-0.16129,-570.01,-1672.5,-83.281,-464.58,-8.9897,-18.572
1547.000000000,-0.16128,-569.19,-1671.7,-83.276,-464.53,-8.9893,-18.570
1548.000000000,-0.16127,-568.50,-1671.1,-83.271,-464.50,-8.9889,-18.569
1549.000000000,-0.16225,1991.2,4114.0,-53.332,-371.11,-9.0237,-20.272
1550.000000000,-0.16202,-571.56,-1673.8,-83.274,-465.75,-9.0154,-18.840
1551.000000000,-0.16174,-570.40,-1672.7,-83.266,-465.26,-9.0074,-18.717
1552.000000000,-0.16155,-569.50,-1671.9,-83.261,-465.06,-9.0013,-18.671
1553.000000000,-0.16333,1990.4,4113.1,-53.322,-372.25,-9.0627,-21.890
1554.000000000,-0.16283,-572.30,-1674.3,-83.263,-466.87,-9.0451,-19.141
1555.000000000,-0.16226,-571.17,-1673.3,-83.255,-466.18,-9.0284,-18.895
1556.000000000,-0.16189,-570.35,-1672.4,-83.251,-465.77,-9.0156,-18.798
1557.000000000,-0.16165,-569.62,-1671.7,-83.248,-465.45,-9.0068,-18.737
1558.000000000,-0.16151,-568.89,-1671.0,-83.244,-465.20,-9.0007,-18.694
1559.000000000,-0.16141,-568.24,-1670.3,-83.239,-465.01,-8.9967,-18.663
1560.000000000,-0.16135,-567.61,-1669.7,-83.235,-464.86,-8.9939,-18.641
1561.000000000,-0.16131,-567.05,-1669.2,-83.232,-464.75,-8.9920,-18.624
1562.000000000,-0.16189,1992.6,4116.3,-53.293,-370.99,-9.0127,-19.666
1563.000000000,-0.16191,1988.8,4111.9,-53.300,-371.52,-9.0133,-19.063
1564.000000000,-0.16189,1985.7,4108.6,-53.303,-371.62,-9.0136,-19.077
1565.000000000,-0.16252,1983.0,4105.8,-53.306,-372.19,-9.0357,-20.186
1566.000000000,-0.16216,-578.49,-1680.0,-83.244,-466.28,-9.0230,-18.912
1567.000000000,-0.16188,1982.6,4105.2,-53.302,-371.52,-9.0154,-18.879
1568.000000000,-0.16194,1979.9,4102.4,-53.308,-371.85,-9.0172,-19.230
1569.000000000,-0.16172,-581.71,-1683.3,-83.247,-465.86,-9.0083,-18.769
1570.000000000,-0.16154,-579.63,-1681.2,-83.240,-465.28,-9.0018,-18.703
1571.000000000,-0.16142,-578.02,-1679.5,-83.236,-465.04,-8.9972,-18.668
1572.000000000,-0.16134,-576.68,-1678.1,-83.232,-464.87,-8.9939,-18.643
1573.000000000,-0.16129,-575.50,-1676.8,-83.229,-464.75,-8.9917,-18.625
1574.000000000,-0.16125,-574.46,-1675.7,-83.225,-464.65,-8.9901,-18.612
1575.000000000,-0.16122,-573.53,-1674.8,-83.221,-464.57,-8.9889,-18.602
1576.000000000,-0.16120,-572.69,-1674.0,-83.218,-464.51,-8.9881,-18.594
1577.000000000,-0.16119,-571.88,-1673.2,-83.215,-464.46,-8.9874,-18.588
1578.000000000,-0.16117,-571.12,-1672.5,-83.212,-464.42,-8.9869,-18.583
1579.000000000,-0.16116,-570.40,-1671.8,-83.209,-464.39,-8.9865,-18.579
1580.000000000,-0.16115,-569.72,-1671.2,-83.206,-464.36,-8.9862,-18.576
1581.000000000,-0.16115,-569.09,-1670.5,-83.202,-464.34,-8.9860,-18.573
1582.000000000,-0.16114,-568.47,-1669.9,-83.199,-464.32,-8.9857,-18.571
1583.000000000,-0.16114,-567.86,-1669.3,-83.196,-464.30,-8.9855,-18.570
1584.000000000,-0.16113,-567.26,-1668.8,-83.192,-464.28,-8.9853,-18.568
1585.000000000,-0.16113,-566.70,-1668.2,-83.188,-464.26,-8.9851,-18.567
1586.000000000,-0.16113,-566.14,-1667.7,-83.184,-464.25,-8.9849,-18.566
1587.000000000,-0.16112,-565.63,-1667.2,-83.180,-464.23,-8.9848,-18.565
1588.000000000,-0.16112,-565.10,-1666.7,-83.177,-464.22,-8.9846,-18.564
1589.000000000,-0.16111,-564.59,-1666.2,-83.173,-464.21,-8.9844,-18.564
1590.000000000,-0.16111,-564.10,-1665.7,-83.169,-464.19,-8.9843,-18.564
1591.000000000,-0.16111,-563.64,-1665.2,-83.165,-464.18,-8.9841,-18.563
1592.000000000,-0.16189,1995.9,4120.1,-53.227,-370.64,-9.0119,-19.908
1593.000000000,-0.16171,-566.96,-1668.2,-83.168,-465.26,-9.0052,-18.777
1594.000000000,-0.16149,-565.88,-1667.3,-83.161,-464.81,-8.9989,-18.681
1595.000000000,-0.16134,-565.03,-1666.5,-83.157,-464.64,-8.9941,-18.644
1596.000000000,-0.16125,-564.32,-1665.9,-83.153,-464.51,-8.9906,-18.621
1597.000000000,-0.16119,-563.70,-1665.3,-83.148,-464.41,-8.9882,-18.605
1598.000000000,-0.16118,1996.0,4120.1,-53.209,-370.19,-8.9883,-18.628
1599.000000000,-0.16115,-566.83,-1668.1,-83.149,-464.69,-8.9863,-18.592
1600.000000000,-0.16112,-565.69,-1667.1,-83.141,-464.31,-8.9853,-18.583
1601.000000000,-0.16264,1994.3,4118.6,-53.201,-371.30,-9.0381,-21.213
1602.000000000,-0.16238,1990.8,4115.0,-53.206,-371.88,-9.0300,-19.168
1603.000000000,-0.16319,1987.9,4111.6,-53.209,-372.72,-9.0606,-21.010
1604.000000000,-0.16261,-573.84,-1674.6,-83.147,-466.77,-9.0407,-19.119
1605.000000000,-0.16210,1986.9,4110.6,-53.205,-371.85,-9.0260,-18.971
1606.000000000,-0.16173,-575.10,-1675.6,-83.147,-465.96,-9.0121,-18.811
1607.000000000,-0.16149,-573.36,-1674.0,-83.140,-465.28,-9.0030,-18.744
1608.000000000,-0.16134,-571.95,-1672.7,-83.135,-464.98,-8.9967,-18.698
1609.000000000,-0.16124,-570.79,-1671.7,-83.131,-464.76,-8.9924,-18.666
1610.000000000,-0.16272,1989.3,4113.5,-53.193,-371.67,-9.0434,-21.292
1611.000000000,-0.16236,1986.0,4109.8,-53.199,-372.12,-9.0313,-19.095
1612.000000000,-0.16693,1983.2,4106.9,-53.203,-375.92,-9.1904,-27.499
1613.000000000,-0.16608,1979.3,4103.7,-53.214,-376.60,-9.1630,-21.147
1614.000000000,-0.16449,1976.2,4100.9,-53.228,-375.82,-9.1168,-19.846
1615.000000000,-0.16362,1973.7,4098.4,-53.244,-375.05,-9.0886,-19.928
1616.000000000,-0.16364,1971.5,4096.4,-53.255,-374.86,-9.0874,-20.712
1617.000000000,-0.16298,1969.5,4094.7,-53.262,-374.27,-9.0630,-19.470
1618.000000000,-0.16235,-591.45,-1690.3,-83.204,-467.72,-9.0394,-19.084
1619.000000000,-0.16193,-589.04,-1687.6,-83.202,-466.70,-9.0230,-18.948
1620.000000000,-0.16166,-587.28,-1685.4,-83.204,-466.15,-9.0117,-18.857
1621.000000000,-0.16149,-585.93,-1683.6,-83.204,-465.75,-9.0041,-18.792
1622.000000000,-0.16138,-584.71,-1681.9,-83.204,-465.44,-8.9989,-18.743
1623.000000000,-0.16130,-583.66,-1680.5,-83.203,-465.21,-8.9952,-18.706
1624.000000000,-0.16124,-582.75,-1679.1,-83.202,-465.02,-8.9927,-18.678
1625.000000000,-0.16120,-581.92,-1677.9,-83.200,-464.88,-8.9909,-18.656
1626.000000000,-0.16117,-581.11,-1676.7,-83.199,-464.77,-8.9896,-18.640
1627.000000000,-0.16115,-580.37,-1675.7,-83.197,-464.68,-8.9887,-18.627
1628.000000000,-0.16114,-579.68,-1674.8,-83.195,-464.62,-8.9882,-18.630
1629.000000000,-0.16112,-579.03,-1674.0,-83.193,-464.56,-8.9876,-18.611
1630.000000000,-0.16111,-578.41,-1673.3,-83.191,-464.51,-8.9871,-18.604
1631.000000000,-0.16110,-577.78,-1672.6,-83.189,-464.47,-8.9867,-18.599
1632.000000000,-0.16109,-577.17,-1671.9,-83.187,-464.44,-8.9864,-18.594
1633.000000000,-0.16108,-576.59,-1671.2,-83.185,-464.42,-8.9861,-18.591
1634.000000000,-0.16107,-576.04,-1670.6,-83.183,-464.39,-8.9859,-18.589
1635.000000000,-0.16107,-575.51,-1670.0,-83.181,-464.37,-8.9857,-18.586
1636.000000000,-0.16108,1984.1,4115.2,-53.244,-370.21,-8.9872,-18.618
1637.000000000,-0.16107,-578.70,-1672.8,-83.189,-464.75,-8.9861,-18.589
1638.000000000,-0.16107,-577.56,-1671.7,-83.185,-464.42,-8.9861,-18.606
1639.000000000,-0.16149,1982.4,4113.3,-53.249,-370.55,-9.0013,-19.313
1640.000000000,-0.16148,1979.0,4109.5,-53.258,-371.03,-9.0010,-18.844
1641.000000000,-0.16134,-583.07,-1676.7,-83.200,-465.18,-8.9960,-18.670
1642.000000000,-0.16124,-581.38,-1675.1,-83.196,-464.73,-8.9925,-18.639
1643.000000000,-0.16117,-580.07,-1673.9,-83.194,-464.60,-8.9899,-18.621
1644.000000000,-0.16114,-578.95,-1672.9,-83.193,-464.51,-8.9883,-18.615
1645.000000000,-0.16111,-577.96,-1672.0,-83.191,-464.44,-8.9870,-18.602
1646.000000000,-0.16109,-577.04,-1671.2,-83.189,-464.39,-8.9861,-18.595
1647.000000000,-0.16113,1982.9,4113.8,-53.252,-370.23,-8.9882,-18.677
1648.000000000,-0.16118,1979.5,4109.9,-53.260,-370.65,-8.9899,-18.713
1649.000000000,-0.16174,1976.6,4106.8,-53.264,-371.16,-9.0092,-19.624
1650.000000000,-0.16232,1974.1,4104.1,-53.268,-371.81,-9.0293,-20.029
1651.000000000,-0.16197,-587.18,-1681.6,-83.207,-465.95,-9.0176,-18.884
1652.000000000,-0.16164,-584.95,-1679.5,-83.200,-465.34,-9.0076,-18.762
1653.000000000,-0.16143,-583.21,-1677.8,-83.197,-465.06,-9.0002,-18.708
1654.000000000,-0.16130,-581.84,-1676.5,-83.193,-464.85,-8.9950,-18.673
1655.000000000,-0.16123,-580.61,-1675.2,-83.191,-464.69,-8.9918,-18.662
1656.000000000,-0.16130,1979.6,4109.1,-53.253,-370.51,-8.9947,-18.846
1657.000000000,-0.16150,1976.4,4105.7,-53.260,-371.04,-9.0015,-19.113
1658.000000000,-0.16180,1973.7,4102.9,-53.263,-371.38,-9.0120,-19.422
1659.000000000,-0.16179,1971.4,4100.4,-53.266,-371.50,-9.0122,-19.110
1660.000000000,-0.16165,1969.4,4098.1,-53.269,-371.45,-9.0079,-18.904
1661.000000000,-0.16152,1967.1,4096.0,-53.271,-371.35,-9.0039,-18.843
1662.000000000,-0.16137,-593.29,-1689.2,-83.209,-465.36,-8.9975,-18.696
1663.000000000,-0.16126,-590.73,-1686.7,-83.201,-464.82,-8.9932,-18.661
1664.000000000,-0.16119,-588.73,-1684.7,-83.197,-464.64,-8.9902,-18.638
1665.000000000,-0.16115,-587.07,-1683.0,-83.193,-464.52,-8.9883,-18.632
1666.000000000,-0.16258,1973.5,4101.7,-53.255,-371.44,-9.0381,-21.137
1667.000000000,-0.16224,-588.53,-1684.6,-83.196,-466.08,-9.0259,-19.026
1668.000000000,-0.16182,-586.70,-1682.8,-83.188,-465.48,-9.0135,-18.822
1669.000000000,-0.16153,-585.31,-1681.4,-83.184,-465.17,-9.0041,-18.748
1670.000000000,-0.16136,-584.01,-1680.1,-83.180,-464.92,-8.9974,-18.702
1671.000000000,-0.16125,-582.84,-1678.9,-83.175,-464.72,-8.9929,-18.670
1672.000000000,-0.16118,-581.74,-1677.8,-83.171,-464.58,-8.9898,-18.646
1673.000000000,-0.16131,1978.4,4106.4,-53.231,-370.44,-8.9948,-18.934
1674.000000000,-0.16132,1975.2,4103.0,-53.237,-370.84,-8.9953,-18.812
1675.000000000,-0.16148,1972.5,4100.1,-53.240,-371.03,-9.0011,-19.090
1676.000000000,-0.16165,1970.2,4097.6,-53.242,-371.23,-9.0068,-19.198
1677.000000000,-0.16146,-591.00,-1687.9,-83.179,-465.32,-9.0000,-18.736
1678.000000000,-0.16133,1970.5,4097.6,-53.236,-370.66,-8.9967,-18.718
1679.000000000,-0.16122,-590.99,-1688.2,-83.177,-465.03,-8.9920,-18.656
1680.000000000,-0.16115,-588.74,-1686.0,-83.169,-464.56,-8.9890,-18.634
1681.000000000,-0.16119,1972.2,4099.0,-53.230,-370.34,-8.9911,-18.776
1682.000000000,-0.16303,1969.5,4096.3,-53.236,-372.16,-9.0542,-21.888
1683.000000000,-0.16256,-591.78,-1689.4,-83.174,-466.49,-9.0377,-19.135
1684.000000000,-0.16202,1969.5,4096.0,-53.232,-371.65,-9.0233,-18.923
1685.000000000,-0.16165,-592.17,-1689.8,-83.174,-465.81,-9.0100,-18.802
1686.000000000,-0.16142,-590.04,-1687.7,-83.166,-465.16,-9.0012,-18.741
1687.000000000,-0.16128,-588.30,-1686.0,-83.162,-464.88,-8.9952,-18.699
1688.000000000,-0.16118,-586.79,-1684.5,-83.159,-464.69,-8.9912,-18.669
1689.000000000,-0.16126,1973.6,4100.0,-53.221,-370.49,-8.9941,-18.880
1690.000000000,-0.16125,1970.5,4096.8,-53.229,-370.83,-8.9936,-18.780
1691.000000000,-0.16117,-591.06,-1689.0,-83.168,-464.96,-8.9899,-18.657
1692.000000000,-0.16111,-588.98,-1687.0,-83.159,-464.50,-8.9877,-18.640
1693.000000000,-0.16106,-587.30,-1685.3,-83.154,-464.37,-8.9859,-18.619
1694.000000000,-0.16103,-585.86,-1683.9,-83.150,-464.28,-8.9845,-18.608
1695.000000000,-0.16101,-584.56,-1682.6,-83.145,-464.21,-8.9835,-18.599
1696.000000000,-0.16099,-583.37,-1681.4,-83.141,-464.16,-8.9829,-18.595
1697.000000000,-0.16144,1976.8,4102.9,-53.201,-370.33,-8.9993,-19.388
1698.000000000,-0.16190,1973.6,4099.6,-53.207,-371.20,-9.0152,-19.690
1699.000000000,-0.16171,1971.0,4096.8,-53.210,-371.28,-9.0098,-18.931
1700.000000000,-0.16180,1968.8,4094.3,-53.213,-371.43,-9.0142,-19.349
1701.000000000,-0.16155,-592.35,-1691.2,-83.150,-465.47,-9.0047,-18.794
1702.000000000,-0.16134,-589.94,-1688.8,-83.142,-464.89,-8.9974,-18.712
1703.000000000,-0.16120,-588.07,-1687.0,-83.137,-464.66,-8.9923,-18.674
1704.000000000,-0.16111,-586.52,-1685.4,-83.132,-464.48,-8.9886,-18.648
1705.000000000,-0.16105,-585.15,-1684.0,-83.128,-464.35,-8.9861,-18.629
1706.000000000,-0.16101,-583.92,-1682.8,-83.124,-464.25,-8.9843,-18.616
1707.000000000,-0.16099,-582.76,-1681.6,-83.120,-464.17,-8.9831,-18.605
1708.000000000,-0.16099,1977.4,4102.7,-53.181,-369.97,-8.9840,-18.636
1709.000000000,-0.16098,-584.97,-1683.9,-83.122,-464.48,-8.9824,-18.598
1710.000000000,-0.16097,-583.41,-1682.4,-83.114,-464.12,-8.9820,-18.607
1711.000000000,-0.16095,-582.12,-1681.1,-83.110,-464.05,-8.9813,-18.588
1712.000000000,-0.16094,-581.00,-1680.0,-83.105,-464.00,-8.9807,-18.583
1713.000000000,-0.16093,-579.99,-1678.9,-83.101,-463.97,-8.9803,-18.580
1714.000000000,-0.16092,-579.06,-1678.0,-83.097,-463.94,-8.9799,-18.577
1715.000000000,-0.16092,-578.17,-1677.1,-83.092,-463.91,-8.9796,-18.575
1716.000000000,-0.16091,-577.32,-1676.2,-83.089,-463.89,-8.9794,-18.573
1717.000000000,-0.16090,-576.50,-1675.5,-83.085,-463.87,-8.9791,-18.572
1718.000000000,-0.16090,-575.71,-1674.9,-83.080,-463.86,-8.9789,-18.571
1719.000000000,-0.16089,-574.96,-1674.2,-83.076,-463.84,-8.9787,-18.570
1720.000000000,-0.16089,-574.20,-1673.6,-83.072,-463.82,-8.9786,-18.569
1721.000000000,-0.16089,-573.47,-1673.0,-83.067,-463.81,-8.9784,-18.568
1722.000000000,-0.16089,-572.75,-1672.4,-83.063,-463.79,-8.9783,-18.567
1723.000000000,-0.16088,-572.05,-1671.8,-83.059,-463.78,-8.9781,-18.566
1724.000000000,-0.16092,1987.7,4113.2,-53.120,-369.64,-8.9802,-18.627
1725.000000000,-0.16090,-574.93,-1674.5,-83.061,-464.18,-8.9790,-18.576
1726.000000000,-0.16089,-573.65,-1673.5,-83.053,-463.84,-8.9785,-18.571
1727.000000000,-0.16091,1986.5,4111.4,-53.113,-369.66,-8.9801,-18.618
1728.000000000,-0.16090,-575.91,-1675.7,-83.054,-464.19,-8.9788,-18.575
1729.000000000,-0.16254,1984.7,4109.0,-53.112,-371.00,-9.0359,-21.411
1730.000000000,-0.16313,1981.6,4105.8,-53.118,-372.29,-9.0570,-20.698
1731.000000000,-0.16577,1979.1,4102.9,-53.122,-374.85,-9.1507,-24.793
1732.000000000,-0.16773,1975.8,4100.0,-53.129,-377.41,-9.2208,-25.420
1733.000000000,-0.16719,1972.5,4097.2,-53.141,-378.09,-9.2086,-22.723
1734.000000000,-0.16559,1969.5,4094.5,-53.158,-377.33,-9.1598,-20.777
1735.000000000,-0.16415,1966.3,4092.0,-53.176,-376.12,-9.1115,-19.922
1736.000000000,-0.16305,-594.17,-1693.2,-83.125,-469.06,-9.0704,-19.380
1737.000000000,-0.16234,-591.87,-1690.6,-83.126,-467.66,-9.0423,-19.166
1738.000000000,-0.16286,1969.1,4094.8,-53.192,-373.43,-9.0574,-20.680
1739.000000000,-0.16252,1966.5,4092.4,-53.206,-373.42,-9.0433,-19.457
1740.000000000,-0.16204,-595.05,-1693.0,-83.151,-467.05,-9.0252,-19.032
1741.000000000,-0.16170,-593.11,-1690.6,-83.149,-466.16,-9.0122,-18.909
1742.000000000,-0.16148,-591.56,-1688.6,-83.149,-465.68,-9.0031,-18.831
1743.000000000,-0.16134,-590.32,-1686.9,-83.148,-465.33,-8.9969,-18.774
1744.000000000,-0.16176,1969.9,4097.9,-53.212,-371.31,-9.0111,-19.604
1745.000000000,-0.16162,1966.6,4094.9,-53.222,-371.57,-9.0057,-18.889
1746.000000000,-0.16143,-595.16,-1690.8,-83.163,-465.57,-8.9987,-18.761
1747.000000000,-0.16130,-593.25,-1688.8,-83.158,-465.00,-8.9938,-18.715
1748.000000000,-0.16122,-591.71,-1687.1,-83.156,-464.80,-8.9905,-18.685
1749.000000000,-0.16117,-590.37,-1685.7,-83.155,-464.64,-8.9881,-18.663
1750.000000000,-0.16114,-589.17,-1684.4,-83.153,-464.53,-8.9867,-18.661
1751.000000000,-0.16111,-588.09,-1683.2,-83.152,-464.44,-8.9854,-18.636
1752.000000000,-0.16109,-587.08,-1682.1,-83.150,-464.37,-8.9845,-18.625
1753.000000000,-0.16108,-586.10,-1681.0,-83.148,-464.31,-8.9838,-18.617
1754.000000000,-0.16107,-585.19,-1680.1,-83.145,-464.26,-8.9833,-18.611
1755.000000000,-0.16106,-584.35,-1679.1,-83.142,-464.23,-8.9829,-18.606
1756.000000000,-0.16105,-583.53,-1678.3,-83.140,-464.19,-8.9826,-18.602
1757.000000000,-0.16104,-582.73,-1677.5,-83.138,-464.17,-8.9823,-18.599
1758.000000000,-0.16104,-581.98,-1676.7,-83.137,-464.14,-8.9821,-18.597
1759.000000000,-0.16104,-581.27,-1676.0,-83.136,-464.12,-8.9819,-18.594
1760.000000000,-0.16104,-580.60,-1675.4,-83.134,-464.11,-8.9817,-18.593
1761.000000000,-0.16104,-579.94,-1674.8,-83.132,-464.09,-8.9816,-18.591
1762.000000000,-0.16103,-579.29,-1674.2,-83.130,-464.08,-8.9815,-18.590
1763.000000000,-0.16103,-578.63,-1673.7,-83.128,-464.06,-8.9813,-18.589
1764.000000000,-0.16103,-577.97,-1673.2,-83.126,-464.05,-8.9812,-18.588
1765.000000000,-0.16103,-577.34,-1672.6,-83.123,-464.04,-8.9811,-18.587
1766.000000000,-0.16104,-576.69,-1672.1,-83.120,-464.03,-8.9813,-18.601
1767.000000000,-0.16104,-576.04,-1671.6,-83.117,-464.02,-8.9811,-18.588
1768.000000000,-0.16103,-575.42,-1671.1,-83.115,-464.01,-8.9810,-18.586
1769.000000000,-0.16103,-574.81,-1670.7,-83.112,-464.00,-8.9808,-18.585
1770.000000000,-0.16103,-574.19,-1670.2,-83.109,-463.98,-8.9807,-18.584
1771.000000000,-0.16102,-573.60,-1669.8,-83.106,-463.97,-8.9806,-18.584
1772.000000000,-0.16102,-573.00,-1669.3,-83.103,-463.96,-8.9805,-18.583
1773.000000000,-0.16102,-572.41,-1668.8,-83.100,-463.95,-8.9803,-18.582
1774.000000000,-0.16104,1987.3,4116.5,-53.161,-369.80,-8.9819,-18.616
1775.000000000,-0.16103,-575.52,-1671.8,-83.104,-464.34,-8.9809,-18.587
1776.000000000,-0.16102,-574.35,-1670.9,-83.097,-464.00,-8.9806,-18.584
1777.000000000,-0.16117,1985.7,4114.4,-53.158,-369.92,-8.9866,-18.844
1778.000000000,-0.16113,-576.84,-1673.3,-83.101,-464.47,-8.9845,-18.624
1779.000000000,-0.16113,1983.6,4111.7,-53.159,-369.97,-8.9856,-18.678
1780.000000000,-0.16109,-578.58,-1675.1,-83.101,-464.46,-8.9834,-18.609
1781.000000000,-0.16106,-576.98,-1673.9,-83.093,-464.08,-8.9821,-18.598
1782.000000000,-0.16104,-575.69,-1672.9,-83.089,-464.01,-8.9812,-18.592
1783.000000000,-0.16102,-574.58,-1672.0,-83.085,-463.96,-8.9806,-18.588
1784.000000000,-0.16101,-573.58,-1671.2,-83.082,-463.92,-8.9800,-18.585
1785.000000000,-0.16100,-572.68,-1670.5,-83.078,-463.89,-8.9796,-18.583
1786.000000000,-0.16099,-571.84,-1669.8,-83.075,-463.87,-8.9793,-18.581
1787.000000000,-0.16098,-571.05,-1669.2,-83.072,-463.85,-8.9791,-18.579
1788.000000000,-0.16097,-570.29,-1668.6,-83.068,-463.83,-8.9788,-18.578
1789.000000000,-0.16097,-569.56,-1668.0,-83.065,-463.81,-8.9786,-18.577
1790.000000000,-0.16096,-568.86,-1667.5,-83.061,-463.79,-8.9784,-18.576
1791.000000000,-0.16096,-568.18,-1667.0,-83.058,-463.78,-8.9782,-18.575
1792.000000000,-0.16095,-567.52,-1666.5,-83.054,-463.76,-8.9781,-18.574
1793.000000000,-0.16095,-566.90,-1666.0,-83.051,-463.75,-8.9779,-18.573
1794.000000000,-0.16094,-566.28,-1665.6,-83.047,-463.74,-8.9777,-18.573
1795.000000000,-0.16094,-565.68,-1665.1,-83.043,-463.72,-8.9776,-18.572
1796.000000000,-0.16093,-565.09,-1664.6,-83.039,-463.71,-8.9774,-18.572
1797.000000000,-0.16093,-564.51,-1664.2,-83.036,-463.70,-8.9772,-18.571
1798.000000000,-0.16092,-563.94,-1663.8,-83.032,-463.69,-8.9771,-18.570
1799.000000000,-0.16092,-563.38,-1663.3,-83.028,-463.67,-8.9769,-18.570
1800.000000000,-0.16091,-562.83,-1662.9,-83.024,-463.66,-8.9767,-18.569
1801.000000000,-0.16135,1996.8,4122.3,-53.085,-369.85,-8.9928,-19.332
1802.000000000,-0.16287,1993.1,4118.9,-53.092,-371.58,-9.0453,-21.481
1803.000000000,-0.16283,1990.0,4115.6,-53.095,-372.09,-9.0454,-19.855
1804.000000000,-0.16220,-571.79,-1671.5,-83.032,-466.02,-9.0259,-18.986
1805.000000000,-0.16173,-570.00,-1670.1,-83.024,-465.25,-9.0105,-18.843
1806.000000000,-0.16143,-568.72,-1669.0,-83.020,-464.86,-8.9996,-18.767
1807.000000000,-0.16124,-567.65,-1668.0,-83.016,-464.56,-8.9921,-18.717
1808.000000000,-0.16113,-566.66,-1667.2,-83.013,-464.33,-8.9871,-18.680
1809.000000000,-0.16105,-565.75,-1666.5,-83.010,-464.16,-8.9837,-18.654
1810.000000000,-0.16100,-564.91,-1665.8,-83.006,-464.03,-8.9814,-18.634
1811.000000000,-0.16104,1995.0,4119.7,-53.067,-369.82,-8.9829,-18.729
1812.000000000,-0.16158,1991.5,4116.3,-53.074,-370.61,-9.0013,-19.616
1813.000000000,-0.16142,-570.56,-1671.2,-83.013,-464.82,-8.9949,-18.768
1814.000000000,-0.16135,1990.2,4114.5,-53.070,-370.25,-8.9943,-18.888
1815.000000000,-0.16121,-571.77,-1672.5,-83.011,-464.63,-8.9886,-18.695
1816.000000000,-0.16110,-570.01,-1671.1,-83.004,-464.15,-8.9845,-18.651
1817.000000000,-0.16102,-568.61,-1670.0,-82.999,-464.00,-8.9815,-18.630
1818.000000000,-0.16099,1991.7,4115.6,-53.060,-369.74,-8.9811,-18.642
1819.000000000,-0.16095,-570.63,-1672.0,-83.001,-464.21,-8.9788,-18.609
1820.000000000,-0.16092,-569.07,-1670.7,-82.993,-463.82,-8.9776,-18.598
1821.000000000,-0.16090,-567.82,-1669.6,-82.989,-463.73,-8.9767,-18.591
1822.000000000,-0.16095,1992.4,4116.0,-53.050,-369.57,-8.9792,-18.695
1823.000000000,-0.16095,1989.2,4112.1,-53.056,-369.96,-8.9796,-18.657
1824.000000000,-0.16092,-572.66,-1674.2,-82.994,-464.14,-8.9777,-18.598
1825.000000000,-0.16090,-570.78,-1672.7,-82.985,-463.75,-8.9769,-18.603
1826.000000000,-0.16087,-569.31,-1671.4,-82.980,-463.67,-8.9760,-18.584
1827.000000000,-0.16086,-568.05,-1670.4,-82.976,-463.62,-8.9752,-18.579
1828.000000000,-0.16086,1992.2,4115.1,-53.037,-369.43,-8.9763,-18.607
1829.000000000,-0.16085,-570.17,-1672.4,-82.978,-463.96,-8.9750,-18.579
1830.000000000,-0.16084,-568.61,-1671.1,-82.970,-463.60,-8.9745,-18.574
1831.000000000,-0.16083,-567.34,-1670.0,-82.966,-463.55,-8.9740,-18.571
1832.000000000,-0.16083,-566.26,-1669.0,-82.961,-463.51,-8.9736,-18.569
1833.000000000,-0.16082,-565.31,-1668.2,-82.957,-463.49,-8.9733,-18.568
1834.000000000,-0.16082,-564.42,-1667.4,-82.952,-463.46,-8.9730,-18.566
1835.000000000,-0.16081,-563.59,-1666.7,-82.948,-463.45,-8.9728,-18.565
1836.000000000,-0.16081,-562.81,-1666.0,-82.943,-463.43,-8.9725,-18.564
1837.000000000,-0.16080,-562.07,-1665.3,-82.939,-463.41,-8.9723,-18.563
1838.000000000,-0.16080,-561.34,-1664.7,-82.934,-463.40,-8.9721,-18.562
1839.000000000,-0.16080,-560.65,-1664.1,-82.929,-463.38,-8.9719,-18.562
1840.000000000,-0.16080,-559.98,-1663.5,-82.925,-463.37,-8.9717,-18.561
1841.000000000,-0.16079,-559.34,-1663.0,-82.920,-463.36,-8.9716,-18.560
1842.000000000,-0.16082,2000.4,4122.4,-52.981,-369.21,-8.9735,-18.614
1843.000000000,-0.16081,-562.38,-1665.7,-82.922,-463.76,-8.9723,-18.569
1844.000000000,-0.16080,-561.17,-1664.7,-82.914,-463.41,-8.9719,-18.564
1845.000000000,-0.16082,1998.9,4121.0,-52.974,-369.23,-8.9734,-18.608
1846.000000000,-0.16083,1995.5,4117.9,-52.980,-369.62,-8.9738,-18.598
1847.000000000,-0.16081,-566.47,-1669.6,-82.918,-463.82,-8.9723,-18.569
1848.000000000,-0.16080,-564.74,-1668.2,-82.909,-463.44,-8.9717,-18.565
1849.000000000,-0.16079,-563.40,-1667.0,-82.904,-463.37,-8.9712,-18.562
1850.000000000,-0.16078,-562.28,-1666.0,-82.899,-463.33,-8.9707,-18.560
1851.000000000,-0.16077,-561.29,-1665.1,-82.895,-463.31,-8.9704,-18.559
1852.000000000,-0.16077,-560.41,-1664.3,-82.891,-463.28,-8.9701,-18.558
1853.000000000,-0.16076,-559.59,-1663.5,-82.886,-463.26,-8.9698,-18.556
1854.000000000,-0.16076,-558.83,-1662.8,-82.881,-463.25,-8.9696,-18.556
1855.000000000,-0.16076,-558.14,-1662.2,-82.877,-463.23,-8.9694,-18.555
1856.000000000,-0.16075,-557.50,-1661.5,-82.872,-463.21,-8.9692,-18.554
1857.000000000,-0.16075,-556.90,-1660.9,-82.867,-463.20,-8.9690,-18.553
1858.000000000,-0.16075,-556.32,-1660.4,-82.863,-463.19,-8.9688,-18.553
1859.000000000,-0.16074,-555.75,-1659.8,-82.858,-463.17,-8.9686,-18.552
1860.000000000,-0.16077,2004.3,4125.5,-52.919,-369.03,-8.9707,-18.612
1861.000000000,-0.16076,-558.61,-1662.6,-82.860,-463.58,-8.9695,-18.562
1862.000000000,-0.16075,-557.48,-1661.7,-82.851,-463.23,-8.9690,-18.557
1863.000000000,-0.16073,-556.57,-1660.8,-82.846,-463.19,-8.9686,-18.554
1864.000000000,-0.16074,2003.7,4124.7,-52.907,-369.01,-8.9698,-18.580
1865.000000000,-0.16073,-559.04,-1663.3,-82.847,-463.55,-8.9686,-18.557
1866.000000000,-0.16072,-557.80,-1662.2,-82.839,-463.20,-8.9682,-18.554
1867.000000000,-0.16071,-556.81,-1661.3,-82.834,-463.15,-8.9678,-18.552
1868.000000000,-0.16070,-555.95,-1660.5,-82.829,-463.12,-8.9675,-18.550
1869.000000000,-0.16069,-555.19,-1659.8,-82.824,-463.10,-8.9672,-18.549
1870.000000000,-0.16080,2005.1,4125.7,-52.885,-369.01,-8.9718,-18.739
1871.000000000,-0.16081,2001.5,4122.5,-52.890,-369.43,-8.9724,-18.644
1872.000000000,-0.16077,-560.58,-1665.1,-82.827,-463.63,-8.9702,-18.576
1873.000000000,-0.16073,-558.95,-1663.7,-82.818,-463.23,-8.9690,-18.565
1874.000000000,-0.16070,-557.72,-1662.6,-82.813,-463.16,-8.9680,-18.559
1875.000000000,-0.16068,-556.69,-1661.6,-82.808,-463.11,-8.9673,-18.556
1876.000000000,-0.16083,2003.7,4124.1,-52.868,-369.04,-8.9734,-18.833
1877.000000000,-0.16126,2000.2,4121.0,-52.874,-369.80,-8.9881,-19.401
1878.000000000,-0.16298,1997.4,4118.4,-52.876,-371.38,-9.0476,-21.931
1879.000000000,-0.16253,1995.0,4115.4,-52.878,-371.60,-9.0338,-19.388
1880.000000000,-0.16188,-566.36,-1670.9,-82.815,-465.42,-9.0139,-18.944
1881.000000000,-0.16147,1994.8,4115.2,-52.871,-370.50,-9.0012,-18.884
1882.000000000,-0.16118,-566.90,-1671.4,-82.813,-464.65,-8.9895,-18.753
1883.000000000,-0.16100,-564.87,-1669.7,-82.805,-464.01,-8.9819,-18.699
1884.000000000,-0.16087,-563.21,-1668.2,-82.800,-463.75,-8.9768,-18.661
1885.000000000,-0.16080,-561.83,-1666.9,-82.796,-463.56,-8.9732,-18.634
1886.000000000,-0.16084,1998.5,4119.0,-52.856,-369.34,-8.9752,-18.782
1887.000000000,-0.16078,-563.77,-1668.6,-82.798,-463.80,-8.9721,-18.626
1888.000000000,-0.16073,-562.15,-1667.2,-82.790,-463.36,-8.9700,-18.601
1889.000000000,-0.16069,-560.82,-1666.1,-82.785,-463.25,-8.9684,-18.588
1890.000000000,-0.16067,-559.66,-1665.0,-82.780,-463.17,-8.9673,-18.578
1891.000000000,-0.16065,-558.68,-1664.1,-82.776,-463.11,-8.9665,-18.570
1892.000000000,-0.16063,-557.82,-1663.2,-82.771,-463.06,-8.9658,-18.564
1893.000000000,-0.16062,-557.01,-1662.4,-82.767,-463.02,-8.9653,-18.560
1894.000000000,-0.16061,-556.25,-1661.6,-82.763,-462.99,-8.9649,-18.556
1895.000000000,-0.16060,-555.53,-1660.9,-82.759,-462.96,-8.9646,-18.553
1896.000000000,-0.16059,-554.85,-1660.2,-82.755,-462.93,-8.9643,-18.551
1897.000000000,-0.16058,-554.21,-1659.6,-82.751,-462.91,-8.9640,-18.549
1898.000000000,-0.16058,-553.58,-1658.9,-82.747,-462.89,-8.9638,-18.548
1899.000000000,-0.16057,-552.98,-1658.3,-82.743,-462.87,-8.9636,-18.546
1900.000000000,-0.16057,-552.40,-1657.7,-82.739,-462.86,-8.9634,-18.545
1901.000000000,-0.16056,-551.84,-1657.1,-82.735,-462.84,-8.9632,-18.544
1902.000000000,-0.16056,-551.28,-1656.6,-82.730,-462.83,-8.9630,-18.543
1903.000000000,-0.16055,-550.75,-1656.0,-82.727,-462.81,-8.9628,-18.542
1904.000000000,-0.16055,-550.27,-1655.5,-82.722,-462.80,-8.9626,-18.542
1905.000000000,-0.16054,-549.79,-1654.9,-82.718,-462.79,-8.9625,-18.541
1906.000000000,-0.16054,-549.32,-1654.4,-82.714,-462.78,-8.9623,-18.541
1907.000000000,-0.16053,-548.87,-1653.9,-82.710,-462.76,-8.9621,-18.540
1908.000000000,-0.16053,-548.42,-1653.4,-82.706,-462.75,-8.9620,-18.539
1909.000000000,-0.16052,-547.98,-1652.9,-82.701,-462.74,-8.9618,-18.539
1910.000000000,-0.16051,-547.55,-1652.5,-82.697,-462.73,-8.9616,-18.538
1911.000000000,-0.16051,-547.14,-1652.0,-82.693,-462.72,-8.9615,-18.538
1912.000000000,-0.16050,-546.73,-1651.5,-82.689,-462.70,-8.9613,-18.537
1913.000000000,-0.16059,2014.1,4133.7,-52.750,-368.61,-8.9653,-18.697
1914.000000000,-0.16057,-549.60,-1654.5,-82.691,-463.16,-8.9638,-18.563
1915.000000000,-0.16053,-548.66,-1653.6,-82.683,-462.81,-8.9628,-18.551
1916.000000000,-0.16051,-547.92,-1652.8,-82.679,-462.75,-8.9620,-18.546
1917.000000000,-0.16050,-547.29,-1652.1,-82.675,-462.72,-8.9615,-18.543
1918.000000000,-0.16048,-546.72,-1651.5,-82.671,-462.69,-8.9610,-18.540
1919.000000000,-0.16047,-546.20,-1651.0,-82.667,-462.67,-8.9606,-18.539
1920.000000000,-0.16047,-545.71,-1650.4,-82.663,-462.64,-8.9603,-18.537
1921.000000000,-0.16046,-545.25,-1649.9,-82.659,-462.63,-8.9601,-18.536
1922.000000000,-0.16045,-544.81,-1649.4,-82.655,-462.61,-8.9599,-18.535
1923.000000000,-0.16045,-544.38,-1648.9,-82.651,-462.59,-8.9597,-18.534
1924.000000000,-0.16044,-543.96,-1648.4,-82.647,-462.58,-8.9595,-18.533
1925.000000000,-0.16044,-543.56,-1647.9,-82.643,-462.57,-8.9593,-18.533
1926.000000000,-0.16043,-543.17,-1647.4,-82.639,-462.55,-8.9591,-18.532
1927.000000000,-0.16042,-542.78,-1647.0,-82.635,-462.54,-8.9589,-18.531
1928.000000000,-0.16042,-542.40,-1646.5,-82.631,-462.53,-8.9588,-18.531
1929.000000000,-0.16041,-542.03,-1646.1,-82.627,-462.51,-8.9586,-18.530
1930.000000000,-0.16046,2019.1,4139.1,-52.689,-368.38,-8.9612,-18.617
1931.000000000,-0.16045,-544.98,-1649.2,-82.630,-462.93,-8.9599,-18.544
1932.000000000,-0.16043,-544.06,-1648.3,-82.623,-462.58,-8.9593,-18.537
1933.000000000,-0.16041,-543.36,-1647.5,-82.619,-462.53,-8.9588,-18.534
1934.000000000,-0.16040,-542.76,-1646.9,-82.615,-462.50,-8.9584,-18.532
1935.000000000,-0.16039,-542.23,-1646.3,-82.611,-462.48,-8.9581,-18.531
1936.000000000,-0.16038,-541.75,-1645.7,-82.608,-462.46,-8.9578,-18.530
1937.000000000,-0.16038,-541.29,-1645.2,-82.604,-462.44,-8.9578,-18.542
1938.000000000,-0.16041,2019.9,4140.1,-52.665,-368.29,-8.9596,-18.582
1939.000000000,-0.16039,-544.14,-1648.1,-82.607,-462.84,-8.9584,-18.537
1940.000000000,-0.16038,-543.20,-1647.2,-82.599,-462.49,-8.9578,-18.532
1941.000000000,-0.16036,-542.46,-1646.4,-82.595,-462.44,-8.9574,-18.530
1942.000000000,-0.16066,2018.9,4139.1,-52.656,-368.50,-8.9687,-19.060
1943.000000000,-0.16059,-544.95,-1649.0,-82.598,-463.06,-8.9654,-18.613
1944.000000000,-0.16049,-543.88,-1648.0,-82.591,-462.67,-8.9626,-18.574
1945.000000000,-0.16043,-543.04,-1647.1,-82.587,-462.57,-8.9605,-18.558
1946.000000000,-0.16039,-542.33,-1646.3,-82.583,-462.50,-8.9589,-18.549
1947.000000000,-0.16036,-541.70,-1645.7,-82.580,-462.44,-8.9579,-18.542
1948.000000000,-0.16034,-541.14,-1645.0,-82.576,-462.40,-8.9571,-18.537
1949.000000000,-0.16042,2020.1,4140.4,-52.637,-368.28,-8.9608,-18.698
1950.000000000,-0.16255,2016.9,4137.1,-52.644,-370.39,-9.0338,-22.260
1951.000000000,-0.16237,2014.0,4134.2,-52.647,-370.90,-9.0287,-19.718
1952.000000000,-0.16167,-548.88,-1653.2,-82.585,-464.79,-9.0078,-18.958
1953.000000000,-0.16117,-547.44,-1651.7,-82.577,-463.99,-8.9915,-18.813
1954.000000000,-0.16086,-546.32,-1650.5,-82.574,-463.57,-8.9799,-18.733
1955.000000000,-0.16066,-545.40,-1649.4,-82.571,-463.26,-8.9720,-18.680
1956.000000000,-0.16054,-544.58,-1648.5,-82.568,-463.02,-8.9667,-18.642
1957.000000000,-0.16045,-543.84,-1647.7,-82.565,-462.84,-8.9631,-18.614
1958.000000000,-0.16040,-543.19,-1646.9,-82.561,-462.70,-8.9607,-18.593
1959.000000000,-0.16036,-542.57,-1646.2,-82.557,-462.59,-8.9589,-18.577
1960.000000000,-0.16033,-541.98,-1645.6,-82.554,-462.50,-8.9577,-18.565
1961.000000000,-0.16031,-541.42,-1645.0,-82.550,-462.43,-8.9568,-18.556
1962.000000000,-0.16030,-540.90,-1644.4,-82.547,-462.38,-8.9561,-18.548
1963.000000000,-0.16029,-540.42,-1643.8,-82.543,-462.33,-8.9556,-18.543
1964.000000000,-0.16029,2020.8,4141.5,-52.604,-368.15,-8.9567,-18.566
1965.000000000,-0.16028,-543.21,-1646.7,-82.547,-462.68,-8.9556,-18.541
1966.000000000,-0.16047,2018.5,4139.1,-52.604,-368.32,-8.9629,-18.878
1967.000000000,-0.16248,2015.6,4136.0,-52.611,-370.34,-9.0321,-22.138
1968.000000000,-0.16201,2012.9,4133.4,-52.615,-370.59,-9.0169,-19.210
1969.000000000,-0.16138,-549.86,-1653.9,-82.553,-464.44,-8.9982,-18.877
1970.000000000,-0.16096,-548.31,-1652.3,-82.546,-463.68,-8.9843,-18.769
1971.000000000,-0.16070,-547.10,-1651.0,-82.543,-463.30,-8.9745,-18.703
1972.000000000,-0.16054,-546.05,-1649.9,-82.540,-463.02,-8.9679,-18.657
1973.000000000,-0.16044,-545.18,-1648.9,-82.537,-462.81,-8.9634,-18.625
1974.000000000,-0.16037,-544.40,-1648.0,-82.534,-462.66,-8.9604,-18.601
1975.000000000,-0.16032,-543.71,-1647.2,-82.531,-462.54,-8.9583,-18.583
1976.000000000,-0.16029,-543.05,-1646.4,-82.529,-462.44,-8.9568,-18.570
1977.000000000,-0.16027,-542.42,-1645.7,-82.526,-462.37,-8.9558,-18.559
1978.000000000,-0.16025,-541.85,-1645.1,-82.523,-462.31,-8.9550,-18.551
1979.000000000,-0.16023,-541.31,-1644.4,-82.520,-462.26,-8.9544,-18.545
1980.000000000,-0.16022,-540.80,-1643.8,-82.517,-462.22,-8.9540,-18.540
1981.000000000,-0.16032,2020.4,4141.5,-52.579,-368.12,-8.9584,-18.724
1982.000000000,-0.16029,-543.52,-1646.6,-82.522,-462.66,-8.9565,-18.564
1983.000000000,-0.16025,-542.52,-1645.6,-82.516,-462.29,-8.9553,-18.548
1984.000000000,-0.16022,-541.72,-1644.7,-82.512,-462.22,-8.9544,-18.540
1985.000000000,-0.16021,-541.04,-1644.0,-82.509,-462.18,-8.9537,-18.535
1986.000000000,-0.16019,-540.42,-1643.3,-82.506,-462.14,-8.9532,-18.532
1987.000000000,-0.16018,-539.85,-1642.6,-82.502,-462.11,-8.9528,-18.529
1988.000000000,-0.16018,-539.32,-1642.0,-82.499,-462.09,-8.9526,-18.535
1989.000000000,-0.16017,-538.82,-1641.4,-82.496,-462.07,-8.9523,-18.526
1990.000000000,-0.16016,-538.34,-1640.8,-82.492,-462.05,-8.9521,-18.524
1991.000000000,-0.16015,-537.89,-1640.3,-82.489,-462.03,-8.9519,-18.524
1992.000000000,-0.16015,-537.46,-1639.8,-82.486,-462.02,-8.9517,-18.522
1993.000000000,-0.16014,-537.06,-1639.3,-82.482,-462.00,-8.9515,-18.521
1994.000000000,-0.16014,-536.67,-1638.8,-82.479,-461.99,-8.9513,-18.520
1995.000000000,-0.16014,-536.31,-1638.3,-82.475,-461.98,-8.9514,-18.534
1996.000000000,-0.16028,2024.8,4146.9,-52.537,-367.93,-8.9571,-18.767
1997.000000000,-0.16024,-539.30,-1641.3,-82.479,-462.48,-8.9551,-18.560
1998.000000000,-0.16019,-538.42,-1640.4,-82.472,-462.12,-8.9537,-18.541
1999.000000000,-0.16019,2023.0,4145.1,-52.533,-367.92,-8.9546,-18.583
2000.000000000,-0.16016,-540.85,-1642.9,-82.476,-462.43,-8.9529,-18.537
2001.000000000,-0.16014,-539.80,-1641.8,-82.469,-462.06,-8.9520,-18.530
2002.000000000,-0.16012,-538.99,-1640.9,-82.465,-462.00,-8.9513,-18.526
2003.000000000,-0.16011,-538.32,-1640.1,-82.461,-461.96,-8.9508,-18.523
2004.000000000,-0.16010,-537.74,-1639.4,-82.457,-461.93,-8.9504,-18.524
2005.000000000,-0.16009,-537.20,-1638.8,-82.454,-461.91,-8.9501,-18.519
2006.000000000,-0.16009,-536.71,-1638.2,-82.450,-461.89,-8.9498,-18.518
2007.000000000,-0.16020,2024.5,4147.2,-52.511,-367.81,-8.9547,-18.724
2008.000000000,-0.16017,-539.46,-1641.0,-82.454,-462.36,-8.9529,-18.549
2009.000000000,-0.16013,-538.48,-1640.0,-82.447,-461.99,-8.9517,-18.533
2010.000000000,-0.16010,-537.70,-1639.2,-82.443,-461.93,-8.9508,-18.527
2011.000000000,-0.16008,-537.04,-1638.4,-82.440,-461.89,-8.9500,-18.523
2012.000000000,-0.16029,2024.3,4147.0,-52.501,-367.87,-8.9580,-18.894
2013.000000000,-0.16061,2021.1,4143.7,-52.508,-368.57,-8.9693,-19.228
2014.000000000,-0.16134,2018.5,4140.9,-52.512,-369.33,-8.9950,-20.170
2015.000000000,-0.16193,2016.1,4138.4,-52.515,-370.09,-9.0161,-20.439
2016.000000000,-0.16177,2014.1,4136.1,-52.518,-370.29,-9.0127,-19.641
2017.000000000,-0.16186,2012.1,4133.9,-52.522,-370.51,-9.0174,-20.024
2018.000000000,-0.16130,-550.55,-1653.0,-82.461,-464.35,-8.9977,-18.952
2019.000000000,-0.16085,-548.66,-1651.0,-82.455,-463.54,-8.9826,-18.802
2020.000000000,-0.16057,-547.23,-1649.5,-82.453,-463.12,-8.9719,-18.724
2021.000000000,-0.16039,-546.02,-1648.1,-82.450,-462.79,-8.9645,-18.671
2022.000000000,-0.16027,-544.98,-1647.0,-82.448,-462.55,-8.9595,-18.633
2023.000000000,-0.16020,-544.03,-1645.9,-82.445,-462.37,-8.9561,-18.605
2024.000000000,-0.16015,-543.20,-1645.0,-82.443,-462.23,-8.9537,-18.584
2025.000000000,-0.16011,-542.45,-1644.1,-82.441,-462.12,-8.9521,-18.568
2026.000000000,-0.16009,-541.77,-1643.3,-82.439,-462.03,-8.9509,-18.556
2027.000000000,-0.16007,-541.11,-1642.6,-82.437,-461.96,-8.9500,-18.547
2028.000000000,-0.16005,-540.48,-1641.9,-82.434,-461.91,-8.9494,-18.539
2029.000000000,-0.16004,-539.88,-1641.2,-82.432,-461.87,-8.9488,-18.534
2030.000000000,-0.16003,-539.32,-1640.5,-82.429,-461.83,-8.9485,-18.529
2031.000000000,-0.16002,-538.79,-1639.9,-82.427,-461.80,-8.9481,-18.525
2032.000000000,-0.16002,-538.27,-1639.3,-82.424,-461.77,-8.9478,-18.522
2033.000000000,-0.16001,-537.77,-1638.7,-82.422,-461.74,-8.9476,-18.520
2034.000000000,-0.16001,-537.29,-1638.2,-82.419,-461.72,-8.9474,-18.518
2035.000000000,-0.16000,-536.83,-1637.6,-82.417,-461.71,-8.9472,-18.517
2036.000000000,-0.16000,-536.37,-1637.1,-82.414,-461.69,-8.9470,-18.515
2037.000000000,-0.16000,-535.93,-1636.6,-82.411,-461.67,-8.9469,-18.514
2038.000000000,-0.16212,2025.2,4148.7,-52.473,-369.20,-9.0205,-22.161
2039.000000000,-0.16171,2022.0,4145.3,-52.480,-369.84,-9.0072,-19.200
2040.000000000,-0.16110,-541.50,-1642.4,-82.419,-463.76,-8.9893,-18.851
2041.000000000,-0.16070,-540.24,-1641.1,-82.412,-463.04,-8.9759,-18.746
2042.000000000,-0.16045,-539.33,-1640.1,-82.409,-462.69,-8.9665,-18.682
2043.000000000,-0.16029,-538.53,-1639.2,-82.406,-462.43,-8.9602,-18.639
2044.000000000,-0.16020,-537.85,-1638.5,-82.403,-462.23,-8.9559,-18.608
2045.000000000,-0.16013,-537.26,-1637.8,-82.400,-462.09,-8.9530,-18.585
2046.000000000,-0.16009,-536.68,-1637.1,-82.397,-461.97,-8.9510,-18.568
2047.000000000,-0.16006,-536.14,-1636.5,-82.393,-461.88,-8.9496,-18.555
2048.000000000,-0.16004,-535.66,-1635.9,-82.390,-461.82,-8.9489,-18.562
2049.000000000,-0.16083,2025.5,4149.4,-52.451,-368.25,-8.9768,-19.926
2050.000000000,-0.16120,2022.2,4146.0,-52.459,-369.13,-8.9898,-19.720
2051.000000000,-0.16159,2019.5,4143.1,-52.463,-369.70,-9.0046,-20.082
2052.000000000,-0.16129,2017.1,4140.5,-52.467,-369.71,-8.9959,-19.209
2053.000000000,-0.16085,-545.80,-1646.7,-82.406,-463.59,-8.9810,-18.807
2054.000000000,-0.16054,-544.23,-1645.0,-82.400,-462.88,-8.9701,-18.717
2055.000000000,-0.16034,-542.99,-1643.7,-82.398,-462.56,-8.9626,-18.663
2056.000000000,-0.16022,-541.94,-1642.5,-82.395,-462.32,-8.9574,-18.626
2057.000000000,-0.16014,-541.05,-1641.5,-82.392,-462.14,-8.9539,-18.599
2058.000000000,-0.16027,2020.5,4144.2,-52.455,-367.99,-8.9586,-18.883
2059.000000000,-0.16053,2017.5,4141.2,-52.463,-368.57,-8.9676,-19.197
2060.000000000,-0.16038,-545.73,-1646.2,-82.402,-462.72,-8.9617,-18.674
2061.000000000,-0.16024,-544.22,-1644.7,-82.396,-462.22,-8.9570,-18.615
2062.000000000,-0.16014,-543.03,-1643.5,-82.393,-462.05,-8.9535,-18.587
2063.000000000,-0.16008,-542.03,-1642.4,-82.390,-461.93,-8.9511,-18.569
2064.000000000,-0.16004,-541.16,-1641.4,-82.388,-461.84,-8.9494,-18.555
2065.000000000,-0.16001,-540.38,-1640.6,-82.385,-461.76,-8.9482,-18.545
2066.000000000,-0.15999,-539.66,-1639.8,-82.383,-461.70,-8.9473,-18.538
2067.000000000,-0.15998,-539.02,-1639.1,-82.380,-461.66,-8.9467,-18.532
2068.000000000,-0.15996,-538.43,-1638.4,-82.378,-461.62,-8.9462,-18.527
2069.000000000,-0.15995,-537.89,-1637.7,-82.375,-461.59,-8.9458,-18.524
