time,DEVILSRIVER
1.000000000000,-18.907
2.000000000000,-18.934
3.000000000000,-18.858
4.000000000000,-18.973
5.000000000000,-18.742
6.000000000000,-18.472
7.000000000000,-18.321
8.000000000000,-18.184
9.000000000000,-19.442
10.00000000000,-19.650
11.00000000000,-17.944
12.00000000000,-17.723
13.00000000000,-17.581
14.00000000000,-17.458
15.00000000000,-17.345
16.00000000000,-17.237
17.00000000000,-17.134
18.00000000000,-17.034
19.00000000000,-16.937
20.00000000000,-16.843
21.00000000000,-16.752
22.00000000000,-16.664
23.00000000000,-16.578
24.00000000000,-16.498
25.00000000000,-16.419
26.00000000000,-16.343
27.00000000000,-16.268
28.00000000000,-16.195
29.00000000000,-16.123
30.00000000000,-16.053
31.00000000000,-15.985
32.00000000000,-15.919
33.00000000000,-15.853
34.00000000000,-15.789
35.00000000000,-15.727
36.00000000000,-15.667
37.00000000000,-15.608
38.00000000000,-15.551
39.00000000000,-15.494
40.00000000000,-15.439
41.00000000000,-15.393
42.00000000000,-15.332
43.00000000000,-15.279
44.00000000000,-15.228
45.00000000000,-15.178
46.00000000000,-15.128
47.00000000000,-15.079
48.00000000000,-15.031
49.00000000000,-14.984
50.00000000000,-14.938
51.00000000000,-14.892
52.00000000000,-14.914
53.00000000000,-14.807
54.00000000000,-14.760
55.00000000000,-14.715
56.00000000000,-14.737
57.00000000000,-14.635
58.00000000000,-14.591
59.00000000000,-14.550
60.00000000000,-14.510
61.00000000000,-14.471
62.00000000000,-14.432
63.00000000000,-14.394
64.00000000000,-14.357
65.00000000000,-14.320
66.00000000000,-14.283
67.00000000000,-14.247
68.00000000000,-14.211
69.00000000000,-14.362
70.00000000000,-14.153
71.00000000000,-14.111
72.00000000000,-14.076
73.00000000000,-14.043
74.00000000000,-14.010
75.00000000000,-13.978
76.00000000000,-13.946
77.00000000000,-13.914
78.00000000000,-13.883
79.00000000000,-13.852
80.00000000000,-13.822
81.00000000000,-13.792
82.00000000000,-13.860
83.00000000000,-13.739
84.00000000000,-13.706
85.00000000000,-13.676
86.00000000000,-13.647
87.00000000000,-13.619
88.00000000000,-13.591
89.00000000000,-13.564
90.00000000000,-13.537
91.00000000000,-13.510
92.00000000000,-13.484
93.00000000000,-13.872
94.00000000000,-13.461
95.00000000000,-13.411
96.00000000000,-13.382
97.00000000000,-13.355
98.00000000000,-13.329
99.00000000000,-13.304
100.0000000000,-13.279
101.0000000000,-13.255
102.0000000000,-13.230
103.0000000000,-13.207
104.0000000000,-13.183
105.0000000000,-13.159
106.0000000000,-13.136
107.0000000000,-13.113
108.0000000000,-13.320
109.0000000000,-13.080
110.0000000000,-13.049
111.0000000000,-13.025
112.0000000000,-13.002
113.0000000000,-12.981
114.0000000000,-12.960
115.0000000000,-12.940
116.0000000000,-12.921
117.0000000000,-12.902
118.0000000000,-13.605
119.0000000000,-14.182
120.0000000000,-12.923
121.0000000000,-12.853
122.0000000000,-13.281
123.0000000000,-12.827
124.0000000000,-12.791
125.0000000000,-12.769
126.0000000000,-12.750
127.0000000000,-12.731
128.0000000000,-12.713
129.0000000000,-12.695
130.0000000000,-12.892
131.0000000000,-12.939
132.0000000000,-12.661
133.0000000000,-12.632
134.0000000000,-12.613
135.0000000000,-12.943
136.0000000000,-12.597
137.0000000000,-12.569
138.0000000000,-12.551
139.0000000000,-12.534
140.0000000000,-12.518
141.0000000000,-12.502
142.0000000000,-12.487
143.0000000000,-12.471
144.0000000000,-13.183
145.0000000000,-12.536
146.0000000000,-13.667
147.0000000000,-12.480
148.0000000000,-12.421
149.0000000000,-12.552
150.0000000000,-12.390
151.0000000000,-12.368
152.0000000000,-12.353
153.0000000000,-12.339
154.0000000000,-12.346
155.0000000000,-12.313
156.0000000000,-12.299
157.0000000000,-12.286
158.0000000000,-12.278
159.0000000000,-12.479
160.0000000000,-12.258
161.0000000000,-12.238
162.0000000000,-12.224
163.0000000000,-12.211
164.0000000000,-12.198
165.0000000000,-12.322
166.0000000000,-13.496
167.0000000000,-12.322
168.0000000000,-12.175
169.0000000000,-12.243
170.0000000000,-12.169
171.0000000000,-12.128
172.0000000000,-12.114
173.0000000000,-12.102
174.0000000000,-12.089
175.0000000000,-12.078
176.0000000000,-12.066
177.0000000000,-12.054
178.0000000000,-12.043
179.0000000000,-12.031
180.0000000000,-12.020
181.0000000000,-12.291
182.0000000000,-12.015
183.0000000000,-12.053
184.0000000000,-11.983
185.0000000000,-11.970
186.0000000000,-11.959
187.0000000000,-11.948
188.0000000000,-11.938
189.0000000000,-11.928
190.0000000000,-11.918
191.0000000000,-11.908
192.0000000000,-11.898
193.0000000000,-11.888
194.0000000000,-11.878
195.0000000000,-11.868
196.0000000000,-11.918
197.0000000000,-12.517
198.0000000000,-12.243
199.0000000000,-11.921
200.0000000000,-11.942
201.0000000000,-11.831
202.0000000000,-11.831
203.0000000000,-11.831
204.0000000000,-11.797
205.0000000000,-11.787
206.0000000000,-11.778
207.0000000000,-11.769
208.0000000000,-11.783
209.0000000000,-11.752
210.0000000000,-11.821
211.0000000000,-11.738
212.0000000000,-11.727
213.0000000000,-11.718
214.0000000000,-11.710
215.0000000000,-11.701
216.0000000000,-11.692
217.0000000000,-11.683
218.0000000000,-11.674
219.0000000000,-11.666
220.0000000000,-11.657
221.0000000000,-11.648
222.0000000000,-11.640
223.0000000000,-11.636
224.0000000000,-11.647
225.0000000000,-11.615
226.0000000000,-11.606
227.0000000000,-11.597
228.0000000000,-11.589
229.0000000000,-11.580
230.0000000000,-11.572
231.0000000000,-11.564
232.0000000000,-11.555
233.0000000000,-11.547
234.0000000000,-11.553
235.0000000000,-11.531
236.0000000000,-11.912
237.0000000000,-11.542
238.0000000000,-11.570
239.0000000000,-12.014
240.0000000000,-11.935
241.0000000000,-11.520
242.0000000000,-11.498
243.0000000000,-11.488
244.0000000000,-11.479
245.0000000000,-11.470
246.0000000000,-11.633
247.0000000000,-11.462
248.0000000000,-11.583
249.0000000000,-11.529
250.0000000000,-11.439
251.0000000000,-11.429
252.0000000000,-11.526
253.0000000000,-11.435
254.0000000000,-11.459
255.0000000000,-11.402
256.0000000000,-11.393
257.0000000000,-11.385
258.0000000000,-11.377
259.0000000000,-11.370
260.0000000000,-11.442
261.0000000000,-11.522
262.0000000000,-11.394
263.0000000000,-12.407
264.0000000000,-12.287
265.0000000000,-11.392
266.0000000000,-11.360
267.0000000000,-11.350
268.0000000000,-11.341
269.0000000000,-11.334
270.0000000000,-11.326
271.0000000000,-11.319
272.0000000000,-11.427
273.0000000000,-11.310
274.0000000000,-11.300
275.0000000000,-11.292
276.0000000000,-11.285
277.0000000000,-11.278
278.0000000000,-11.271
279.0000000000,-11.265
280.0000000000,-11.257
281.0000000000,-11.250
282.0000000000,-11.243
283.0000000000,-11.236
284.0000000000,-11.229
285.0000000000,-11.222
286.0000000000,-11.217
287.0000000000,-11.300
288.0000000000,-11.374
289.0000000000,-11.762
290.0000000000,-11.233
291.0000000000,-11.201
292.0000000000,-11.195
293.0000000000,-11.186
294.0000000000,-11.179
295.0000000000,-11.172
296.0000000000,-11.166
297.0000000000,-11.159
298.0000000000,-11.152
299.0000000000,-11.146
300.0000000000,-11.139
301.0000000000,-11.133
302.0000000000,-11.126
303.0000000000,-11.119
304.0000000000,-11.116
305.0000000000,-11.107
306.0000000000,-11.100
307.0000000000,-11.094
308.0000000000,-11.137
309.0000000000,-11.097
310.0000000000,-11.119
311.0000000000,-11.107
312.0000000000,-11.067
313.0000000000,-11.099
314.0000000000,-11.056
315.0000000000,-11.049
316.0000000000,-11.049
317.0000000000,-11.038
318.0000000000,-11.030
319.0000000000,-11.024
320.0000000000,-11.017
321.0000000000,-11.011
322.0000000000,-11.005
323.0000000000,-10.999
324.0000000000,-10.992
325.0000000000,-10.986
326.0000000000,-10.992
327.0000000000,-10.986
328.0000000000,-11.055
329.0000000000,-11.041
330.0000000000,-10.965
331.0000000000,-10.957
332.0000000000,-10.950
333.0000000000,-10.944
334.0000000000,-10.938
335.0000000000,-10.932
336.0000000000,-10.926
337.0000000000,-10.919
338.0000000000,-10.913
339.0000000000,-10.907
340.0000000000,-10.916
341.0000000000,-10.896
342.0000000000,-10.890
343.0000000000,-10.884
344.0000000000,-10.878
345.0000000000,-10.872
346.0000000000,-10.866
347.0000000000,-10.860
348.0000000000,-10.854
349.0000000000,-10.848
350.0000000000,-10.842
351.0000000000,-10.836
352.0000000000,-10.830
353.0000000000,-10.824
354.0000000000,-10.818
355.0000000000,-10.859
356.0000000000,-10.828
357.0000000000,-10.804
358.0000000000,-10.798
359.0000000000,-10.792
360.0000000000,-10.802
361.0000000000,-10.813
362.0000000000,-10.805
363.0000000000,-10.773
364.0000000000,-10.767
365.0000000000,-10.761
366.0000000000,-10.755
367.0000000000,-10.749
368.0000000000,-10.744
369.0000000000,-10.738
370.0000000000,-10.732
371.0000000000,-10.726
372.0000000000,-10.721
373.0000000000,-10.715
374.0000000000,-10.709
375.0000000000,-10.704
376.0000000000,-10.698
377.0000000000,-10.692
378.0000000000,-10.687
379.0000000000,-10.681
380.0000000000,-10.675
381.0000000000,-10.670
382.0000000000,-10.664
383.0000000000,-10.658
384.0000000000,-10.653
385.0000000000,-10.647
386.0000000000,-10.642
387.0000000000,-10.636
388.0000000000,-10.630
389.0000000000,-10.628
390.0000000000,-10.620
391.0000000000,-10.614
392.0000000000,-10.608
393.0000000000,-10.603
394.0000000000,-10.597
395.0000000000,-10.592
396.0000000000,-10.586
397.0000000000,-10.581
398.0000000000,-10.575
399.0000000000,-10.570
400.0000000000,-10.564
401.0000000000,-10.558
402.0000000000,-10.553
403.0000000000,-10.547
404.0000000000,-10.542
405.0000000000,-10.536
406.0000000000,-10.531
407.0000000000,-10.525
408.0000000000,-10.519
409.0000000000,-10.514
410.0000000000,-10.508
411.0000000000,-10.503
412.0000000000,-10.497
413.0000000000,-10.492
414.0000000000,-10.486
415.0000000000,-10.481
416.0000000000,-10.475
417.0000000000,-10.470
418.0000000000,-10.464
419.0000000000,-10.459
420.0000000000,-10.454
421.0000000000,-10.450
422.0000000000,-10.466
423.0000000000,-10.447
424.0000000000,-10.435
425.0000000000,-10.429
426.0000000000,-10.425
427.0000000000,-10.419
428.0000000000,-10.413
429.0000000000,-10.408
430.0000000000,-10.403
431.0000000000,-10.397
432.0000000000,-10.392
433.0000000000,-10.387
434.0000000000,-10.382
435.0000000000,-10.376
436.0000000000,-10.371
437.0000000000,-10.365
438.0000000000,-10.360
439.0000000000,-10.355
440.0000000000,-10.349
441.0000000000,-10.344
442.0000000000,-10.339
443.0000000000,-10.333
444.0000000000,-10.328
445.0000000000,-10.323
446.0000000000,-10.318
447.0000000000,-10.312
448.0000000000,-10.311
449.0000000000,-10.302
450.0000000000,-10.297
451.0000000000,-10.292
452.0000000000,-10.287
453.0000000000,-10.281
454.0000000000,-10.276
455.0000000000,-10.271
456.0000000000,-10.266
457.0000000000,-10.260
458.0000000000,-10.255
459.0000000000,-10.264
460.0000000000,-10.247
461.0000000000,-10.242
462.0000000000,-10.236
463.0000000000,-10.232
464.0000000000,-10.226
465.0000000000,-10.221
466.0000000000,-10.216
467.0000000000,-10.210
468.0000000000,-10.205
469.0000000000,-10.200
470.0000000000,-10.195
471.0000000000,-10.190
472.0000000000,-10.185
473.0000000000,-10.180
474.0000000000,-10.174
475.0000000000,-10.171
476.0000000000,-10.164
477.0000000000,-10.159
478.0000000000,-10.154
479.0000000000,-10.149
480.0000000000,-10.144
481.0000000000,-10.139
482.0000000000,-10.134
483.0000000000,-10.129
484.0000000000,-10.124
485.0000000000,-10.118
486.0000000000,-10.113
487.0000000000,-10.108
488.0000000000,-10.103
489.0000000000,-10.098
490.0000000000,-10.093
491.0000000000,-10.088
492.0000000000,-10.091
493.0000000000,-10.080
494.0000000000,-10.078
495.0000000000,-10.077
496.0000000000,-10.066
497.0000000000,-10.061
498.0000000000,-10.064
499.0000000000,-10.054
500.0000000000,-10.048
501.0000000000,-10.043
502.0000000000,-10.038
503.0000000000,-10.033
504.0000000000,-10.028
505.0000000000,-10.023
506.0000000000,-10.018
507.0000000000,-10.013
508.0000000000,-10.010
509.0000000000,-10.003
510.0000000000,-10.005
511.0000000000,-10.043
512.0000000000,-10.002
513.0000000000,-9.9940
514.0000000000,-9.9890
515.0000000000,-9.9840
516.0000000000,-9.9790
517.0000000000,-9.9741
518.0000000000,-9.9691
519.0000000000,-9.9642
520.0000000000,-9.9592
521.0000000000,-9.9543
522.0000000000,-9.9493
523.0000000000,-9.9444
524.0000000000,-9.9395
525.0000000000,-9.9351
526.0000000000,-9.9302
527.0000000000,-9.9249
528.0000000000,-9.9212
529.0000000000,-9.9236
530.0000000000,-9.9277
531.0000000000,-9.9110
532.0000000000,-9.9059
533.0000000000,-9.9011
534.0000000000,-9.8962
535.0000000000,-9.8913
536.0000000000,-9.9778
537.0000000000,-9.9452
538.0000000000,-9.9178
539.0000000000,-9.9014
540.0000000000,-9.8969
541.0000000000,-9.9263
542.0000000000,-9.8939
543.0000000000,-9.8888
544.0000000000,-9.8842
545.0000000000,-9.8791
546.0000000000,-9.8742
547.0000000000,-9.8693
548.0000000000,-9.8644
549.0000000000,-9.8596
550.0000000000,-9.8547
551.0000000000,-9.8498
552.0000000000,-9.8449
553.0000000000,-9.8401
554.0000000000,-9.8352
555.0000000000,-9.8304
556.0000000000,-9.8258
557.0000000000,-9.8211
558.0000000000,-9.8206
559.0000000000,-9.8127
560.0000000000,-9.8078
561.0000000000,-9.8029
562.0000000000,-9.8041
563.0000000000,-9.8025
564.0000000000,-9.7981
565.0000000000,-9.7895
566.0000000000,-9.7847
567.0000000000,-9.7798
568.0000000000,-9.7750
569.0000000000,-9.7702
570.0000000000,-9.7654
571.0000000000,-9.7632
572.0000000000,-9.7566
573.0000000000,-9.7518
574.0000000000,-9.7470
575.0000000000,-9.7422
576.0000000000,-9.7374
577.0000000000,-9.7327
578.0000000000,-9.7279
579.0000000000,-9.7339
580.0000000000,-9.7497
581.0000000000,-9.7261
582.0000000000,-9.7210
583.0000000000,-9.7163
584.0000000000,-9.7115
585.0000000000,-9.7068
586.0000000000,-9.7021
587.0000000000,-9.6974
588.0000000000,-9.6927
589.0000000000,-9.6897
590.0000000000,-9.6907
591.0000000000,-9.6817
592.0000000000,-9.6769
593.0000000000,-9.6722
594.0000000000,-9.6686
595.0000000000,-9.6704
596.0000000000,-9.6715
597.0000000000,-9.6601
598.0000000000,-9.6554
599.0000000000,-9.6507
600.0000000000,-9.6460
601.0000000000,-9.6413
602.0000000000,-9.6367
603.0000000000,-9.6320
604.0000000000,-9.6274
605.0000000000,-9.6229
606.0000000000,-9.6182
607.0000000000,-9.6141
608.0000000000,-9.6096
609.0000000000,-9.6050
610.0000000000,-9.6004
611.0000000000,-9.5958
612.0000000000,-9.5913
613.0000000000,-9.5904
614.0000000000,-9.5859
615.0000000000,-9.5810
616.0000000000,-9.5794
617.0000000000,-9.5738
618.0000000000,-9.5692
619.0000000000,-9.5647
620.0000000000,-9.5602
621.0000000000,-9.5564
622.0000000000,-9.5525
623.0000000000,-9.5480
624.0000000000,-9.5435
625.0000000000,-9.5394
626.0000000000,-9.5348
627.0000000000,-9.5350
628.0000000000,-9.5309
629.0000000000,-9.5286
630.0000000000,-9.5258
631.0000000000,-9.5209
632.0000000000,-9.5164
633.0000000000,-9.5120
634.0000000000,-9.5076
635.0000000000,-9.5181
636.0000000000,-9.5112
637.0000000000,-9.5060
638.0000000000,-9.5015
639.0000000000,-9.4970
640.0000000000,-9.4924
641.0000000000,-9.4879
642.0000000000,-9.4834
643.0000000000,-9.4789
644.0000000000,-9.4745
645.0000000000,-9.4700
646.0000000000,-9.4655
647.0000000000,-9.4610
648.0000000000,-9.4565
649.0000000000,-9.4563
650.0000000000,-9.4518
651.0000000000,-9.4474
652.0000000000,-9.4429
653.0000000000,-9.4385
654.0000000000,-9.4340
655.0000000000,-9.4296
656.0000000000,-9.4251
657.0000000000,-9.4207
658.0000000000,-9.4163
659.0000000000,-9.4120
660.0000000000,-9.4084
661.0000000000,-9.4064
662.0000000000,-9.4020
663.0000000000,-9.3975
664.0000000000,-9.3931
665.0000000000,-9.3887
666.0000000000,-9.3843
667.0000000000,-9.3799
668.0000000000,-9.3755
669.0000000000,-9.3712
670.0000000000,-9.3668
671.0000000000,-9.3624
672.0000000000,-9.3580
673.0000000000,-9.3537
674.0000000000,-9.3636
675.0000000000,-9.3671
676.0000000000,-9.3629
677.0000000000,-9.3587
678.0000000000,-9.3543
679.0000000000,-9.3500
680.0000000000,-9.3456
681.0000000000,-9.3412
682.0000000000,-9.3369
683.0000000000,-9.3325
684.0000000000,-9.3281
685.0000000000,-9.3238
686.0000000000,-9.3195
687.0000000000,-9.3151
688.0000000000,-9.3108
689.0000000000,-9.3065
690.0000000000,-9.3021
691.0000000000,-9.2978
692.0000000000,-9.2948
693.0000000000,-9.2905
694.0000000000,-9.2862
695.0000000000,-9.2819
696.0000000000,-9.2776
697.0000000000,-9.2733
698.0000000000,-9.2690
699.0000000000,-9.2647
700.0000000000,-9.2605
701.0000000000,-9.2562
702.0000000000,-9.2519
703.0000000000,-9.2477
704.0000000000,-9.2434
705.0000000000,-9.2392
706.0000000000,-9.2349
707.0000000000,-9.2307
708.0000000000,-9.2265
709.0000000000,-9.2223
710.0000000000,-9.2181
711.0000000000,-9.2139
712.0000000000,-9.2097
713.0000000000,-9.2055
714.0000000000,-9.2013
715.0000000000,-9.1971
716.0000000000,-9.1929
717.0000000000,-9.1887
718.0000000000,-9.1847
719.0000000000,-9.1805
720.0000000000,-9.1763
721.0000000000,-9.1722
722.0000000000,-9.1681
723.0000000000,-9.1642
724.0000000000,-9.1600
725.0000000000,-9.1559
726.0000000000,-9.1517
727.0000000000,-9.1531
728.0000000000,-9.1492
729.0000000000,-9.1451
730.0000000000,-9.1412
731.0000000000,-9.1382
732.0000000000,-9.1357
733.0000000000,-9.1335
734.0000000000,-9.1294
735.0000000000,-9.1252
736.0000000000,-9.1211
737.0000000000,-9.1170
738.0000000000,-9.1129
739.0000000000,-9.1090
740.0000000000,-9.1075
741.0000000000,-9.1037
742.0000000000,-9.0996
743.0000000000,-9.0956
744.0000000000,-9.0915
745.0000000000,-9.0874
746.0000000000,-9.0833
747.0000000000,-9.0793
748.0000000000,-9.0752
749.0000000000,-9.0712
750.0000000000,-9.0671
751.0000000000,-9.0631
752.0000000000,-9.0608
753.0000000000,-9.0588
754.0000000000,-9.0549
755.0000000000,-9.0509
756.0000000000,-9.0469
757.0000000000,-9.0429
758.0000000000,-9.0389
759.0000000000,-9.0349
760.0000000000,-9.0309
761.0000000000,-9.0285
762.0000000000,-9.0267
763.0000000000,-9.0227
764.0000000000,-9.0187
765.0000000000,-9.0149
766.0000000000,-9.0109
767.0000000000,-9.0069
768.0000000000,-9.0029
769.0000000000,-8.9990
770.0000000000,-8.9950
771.0000000000,-8.9911
772.0000000000,-8.9871
773.0000000000,-8.9832
774.0000000000,-8.9793
775.0000000000,-8.9753
776.0000000000,-8.9714
777.0000000000,-8.9675
778.0000000000,-8.9638
779.0000000000,-8.9599
780.0000000000,-8.9560
781.0000000000,-8.9521
782.0000000000,-8.9482
783.0000000000,-8.9443
784.0000000000,-8.9404
785.0000000000,-8.9365
786.0000000000,-8.9327
787.0000000000,-8.9288
788.0000000000,-8.9249
789.0000000000,-8.9217
790.0000000000,-8.9181
791.0000000000,-8.9143
792.0000000000,-8.9104
793.0000000000,-8.9066
794.0000000000,-8.9052
795.0000000000,-8.9014
796.0000000000,-8.8975
797.0000000000,-8.8945
798.0000000000,-8.8909
799.0000000000,-8.8874
800.0000000000,-8.8836
801.0000000000,-8.8798
802.0000000000,-8.8760
803.0000000000,-8.8722
804.0000000000,-8.8684
805.0000000000,-8.8646
806.0000000000,-8.8608
807.0000000000,-8.8575
808.0000000000,-8.8538
809.0000000000,-8.8528
810.0000000000,-8.8589
811.0000000000,-8.8608
812.0000000000,-8.8570
813.0000000000,-8.8532
814.0000000000,-8.8494
815.0000000000,-8.8460
816.0000000000,-8.8422
817.0000000000,-8.8385
818.0000000000,-8.8347
819.0000000000,-8.8310
820.0000000000,-8.8272
821.0000000000,-8.8235
822.0000000000,-8.8197
823.0000000000,-8.8160
824.0000000000,-8.8123
825.0000000000,-8.8085
826.0000000000,-8.8053
827.0000000000,-8.8016
828.0000000000,-8.7980
829.0000000000,-8.7955
830.0000000000,-8.7918
831.0000000000,-8.7881
832.0000000000,-8.7852
833.0000000000,-8.7858
834.0000000000,-8.7821
835.0000000000,-8.7784
836.0000000000,-8.7770
837.0000000000,-8.7739
838.0000000000,-8.7736
839.0000000000,-8.7700
840.0000000000,-8.7663
841.0000000000,-8.7626
842.0000000000,-8.7590
843.0000000000,-8.7553
844.0000000000,-8.7541
845.0000000000,-8.7505
846.0000000000,-8.7468
847.0000000000,-8.7473
848.0000000000,-8.7436
849.0000000000,-8.7400
850.0000000000,-8.7364
851.0000000000,-8.7327
852.0000000000,-8.7291
853.0000000000,-8.7255
854.0000000000,-8.7218
855.0000000000,-8.7183
856.0000000000,-8.7147
857.0000000000,-8.7112
858.0000000000,-8.7076
859.0000000000,-8.7040
860.0000000000,-8.7004
861.0000000000,-8.7096
862.0000000000,-8.7154
863.0000000000,-8.7188
864.0000000000,-8.7178
865.0000000000,-8.7155
866.0000000000,-8.7172
867.0000000000,-8.7231
868.0000000000,-8.7195
869.0000000000,-8.7159
870.0000000000,-8.7122
871.0000000000,-8.7128
872.0000000000,-8.7100
873.0000000000,-8.7066
874.0000000000,-8.7054
875.0000000000,-8.7020
876.0000000000,-8.6994
877.0000000000,-8.6958
878.0000000000,-8.6922
879.0000000000,-8.6993
880.0000000000,-8.6959
881.0000000000,-8.7006
882.0000000000,-8.6970
883.0000000000,-8.6933
884.0000000000,-8.6897
885.0000000000,-8.6861
886.0000000000,-8.6825
887.0000000000,-8.6789
888.0000000000,-8.6753
889.0000000000,-8.6717
890.0000000000,-8.6681
891.0000000000,-8.6645
892.0000000000,-8.6609
893.0000000000,-8.6573
894.0000000000,-8.6547
895.0000000000,-8.6582
896.0000000000,-8.6554
897.0000000000,-8.6552
898.0000000000,-8.6530
899.0000000000,-8.6496
900.0000000000,-8.6461
901.0000000000,-8.6459
902.0000000000,-8.6426
903.0000000000,-8.6391
904.0000000000,-8.6363
905.0000000000,-8.6328
906.0000000000,-8.6293
907.0000000000,-8.6257
908.0000000000,-8.6264
909.0000000000,-8.6267
910.0000000000,-8.6234
911.0000000000,-8.6199
912.0000000000,-8.6173
913.0000000000,-8.6138
914.0000000000,-8.6103
915.0000000000,-8.6067
916.0000000000,-8.6032
917.0000000000,-8.5997
918.0000000000,-8.5962
919.0000000000,-8.5970
920.0000000000,-8.5935
921.0000000000,-8.5900
922.0000000000,-8.5865
923.0000000000,-8.5831
924.0000000000,-8.5796
925.0000000000,-8.5761
926.0000000000,-8.5726
927.0000000000,-8.5692
928.0000000000,-8.5657
929.0000000000,-8.5622
930.0000000000,-8.5588
931.0000000000,-8.5553
932.0000000000,-8.5519
933.0000000000,-8.5484
934.0000000000,-8.5450
935.0000000000,-8.5416
936.0000000000,-8.5382
937.0000000000,-8.5347
938.0000000000,-8.5313
939.0000000000,-8.5279
940.0000000000,-8.5245
941.0000000000,-8.5211
942.0000000000,-8.5177
943.0000000000,-8.5155
944.0000000000,-8.5134
945.0000000000,-8.5100
946.0000000000,-8.5066
947.0000000000,-8.5032
948.0000000000,-8.4999
949.0000000000,-8.4965
950.0000000000,-8.4931
951.0000000000,-8.4898
952.0000000000,-8.4864
953.0000000000,-8.4831
954.0000000000,-8.4797
955.0000000000,-8.4776
956.0000000000,-8.4752
957.0000000000,-8.4737
958.0000000000,-8.4730
959.0000000000,-8.4697
960.0000000000,-8.4663
961.0000000000,-8.4630
962.0000000000,-8.4633
963.0000000000,-8.4616
964.0000000000,-8.4583
965.0000000000,-8.4550
966.0000000000,-8.4517
967.0000000000,-8.4484
968.0000000000,-8.4458
969.0000000000,-8.4434
970.0000000000,-8.4401
971.0000000000,-8.4368
972.0000000000,-8.4335
973.0000000000,-8.4307
974.0000000000,-8.4275
975.0000000000,-8.4242
976.0000000000,-8.4209
977.0000000000,-8.4177
978.0000000000,-8.4144
979.0000000000,-8.4112
980.0000000000,-8.4079
981.0000000000,-8.4047
982.0000000000,-8.4015
983.0000000000,-8.4004
984.0000000000,-8.3971
985.0000000000,-8.3951
986.0000000000,-8.3919
987.0000000000,-8.3887
988.0000000000,-8.3855
989.0000000000,-8.3823
990.0000000000,-8.3791
991.0000000000,-8.3759
992.0000000000,-8.3727
993.0000000000,-8.3695
994.0000000000,-8.3663
995.0000000000,-8.3632
996.0000000000,-8.3600
997.0000000000,-8.3568
998.0000000000,-8.3537
999.0000000000,-8.3505
1000.000000000,-8.3482
1001.000000000,-8.3451
1002.000000000,-8.3419
1003.000000000,-8.3388
1004.000000000,-8.3356
1005.000000000,-8.3325
1006.000000000,-8.3294
1007.000000000,-8.3263
1008.000000000,-8.3231
1009.000000000,-8.3200
1010.000000000,-8.3169
1011.000000000,-8.3138
1012.000000000,-8.3206
1013.000000000,-8.3191
1014.000000000,-8.3160
1015.000000000,-8.3129
1016.000000000,-8.3097
1017.000000000,-8.3066
1018.000000000,-8.3035
1019.000000000,-8.3005
1020.000000000,-8.2974
1021.000000000,-8.2943
1022.000000000,-8.2912
1023.000000000,-8.2881
1024.000000000,-8.2851
1025.000000000,-8.2826
1026.000000000,-8.2806
1027.000000000,-8.2981
1028.000000000,-8.3040
1029.000000000,-8.3009
1030.000000000,-8.2978
1031.000000000,-8.2947
1032.000000000,-8.2916
1033.000000000,-8.2893
1034.000000000,-8.2982
1035.000000000,-8.2951
1036.000000000,-8.2920
1037.000000000,-8.2889
1038.000000000,-8.2858
1039.000000000,-8.2827
1040.000000000,-8.2796
1041.000000000,-8.2771
1042.000000000,-8.2745
1043.000000000,-8.2714
1044.000000000,-8.2683
1045.000000000,-8.2652
1046.000000000,-8.2622
1047.000000000,-8.2591
1048.000000000,-8.2563
1049.000000000,-8.2541
1050.000000000,-8.2513
1051.000000000,-8.2485
1052.000000000,-8.2455
1053.000000000,-8.2424
1054.000000000,-8.2394
1055.000000000,-8.2364
1056.000000000,-8.2334
1057.000000000,-8.2304
1058.000000000,-8.2273
1059.000000000,-8.2243
1060.000000000,-8.2217
1061.000000000,-8.2205
1062.000000000,-8.2249
1063.000000000,-8.2223
1064.000000000,-8.2193
1065.000000000,-8.2163
1066.000000000,-8.2133
1067.000000000,-8.2103
1068.000000000,-8.2073
1069.000000000,-8.2043
1070.000000000,-8.2013
1071.000000000,-8.1984
1072.000000000,-8.1954
1073.000000000,-8.1924
1074.000000000,-8.1895
1075.000000000,-8.1865
1076.000000000,-8.1836
1077.000000000,-8.1894
1078.000000000,-8.1864
1079.000000000,-8.1835
1080.000000000,-8.1805
1081.000000000,-8.1776
1082.000000000,-8.1746
1083.000000000,-8.1717
1084.000000000,-8.1688
1085.000000000,-8.1658
1086.000000000,-8.1629
1087.000000000,-8.1600
1088.000000000,-8.1571
1089.000000000,-8.1542
1090.000000000,-8.1513
1091.000000000,-8.1558
1092.000000000,-8.1544
1093.000000000,-8.1515
1094.000000000,-8.1486
1095.000000000,-8.1457
1096.000000000,-8.1428
1097.000000000,-8.1400
1098.000000000,-8.1384
1099.000000000,-8.1356
1100.000000000,-8.1327
1101.000000000,-8.1298
1102.000000000,-8.1269
1103.000000000,-8.1240
1104.000000000,-8.1212
1105.000000000,-8.1183
1106.000000000,-8.1155
1107.000000000,-8.1126
1108.000000000,-8.1098
1109.000000000,-8.1069
1110.000000000,-8.1041
1111.000000000,-8.1012
1112.000000000,-8.0984
1113.000000000,-8.0956
1114.000000000,-8.0928
1115.000000000,-8.0899
1116.000000000,-8.0871
1117.000000000,-8.0843
1118.000000000,-8.0815
1119.000000000,-8.0787
1120.000000000,-8.0759
1121.000000000,-8.0731
1122.000000000,-8.0749
1123.000000000,-8.0721
1124.000000000,-8.0693
1125.000000000,-8.0665
1126.000000000,-8.0637
1127.000000000,-8.0609
1128.000000000,-8.0582
1129.000000000,-8.0554
1130.000000000,-8.0526
1131.000000000,-8.0499
1132.000000000,-8.0471
1133.000000000,-8.0444
1134.000000000,-8.0416
1135.000000000,-8.0389
1136.000000000,-8.0361
1137.000000000,-8.0334
1138.000000000,-8.0307
1139.000000000,-8.0279
1140.000000000,-8.0252
1141.000000000,-8.0225
1142.000000000,-8.0198
1143.000000000,-8.0171
1144.000000000,-8.0144
1145.000000000,-8.0117
1146.000000000,-8.0090
1147.000000000,-8.0063
1148.000000000,-8.0053
1149.000000000,-8.0074
1150.000000000,-8.0047
1151.000000000,-8.0020
1152.000000000,-7.9993
1153.000000000,-7.9966
1154.000000000,-7.9939
1155.000000000,-7.9913
1156.000000000,-7.9886
1157.000000000,-7.9859
1158.000000000,-7.9833
1159.000000000,-7.9806
1160.000000000,-7.9779
1161.000000000,-7.9753
1162.000000000,-7.9726
1163.000000000,-7.9780
1164.000000000,-7.9804
1165.000000000,-7.9853
1166.000000000,-7.9901
1167.000000000,-7.9920
1168.000000000,-7.9893
1169.000000000,-7.9866
1170.000000000,-7.9839
1171.000000000,-7.9812
1172.000000000,-7.9787
1173.000000000,-7.9760
1174.000000000,-7.9770
1175.000000000,-7.9744
1176.000000000,-7.9717
1177.000000000,-7.9690
1178.000000000,-7.9664
1179.000000000,-7.9642
1180.000000000,-7.9616
1181.000000000,-7.9589
1182.000000000,-7.9563
1183.000000000,-7.9536
1184.000000000,-7.9510
1185.000000000,-7.9484
1186.000000000,-7.9457
1187.000000000,-7.9432
1188.000000000,-7.9406
1189.000000000,-7.9380
1190.000000000,-7.9353
1191.000000000,-7.9327
1192.000000000,-7.9301
1193.000000000,-7.9275
1194.000000000,-7.9249
1195.000000000,-7.9223
1196.000000000,-7.9198
1197.000000000,-7.9173
1198.000000000,-7.9147
1199.000000000,-7.9154
1200.000000000,-7.9129
1201.000000000,-7.9103
1202.000000000,-7.9077
1203.000000000,-7.9270
1204.000000000,-7.9292
1205.000000000,-7.9267
1206.000000000,-7.9242
1207.000000000,-7.9216
1208.000000000,-7.9191
1209.000000000,-7.9165
1210.000000000,-7.9142
1211.000000000,-7.9117
1212.000000000,-7.9091
1213.000000000,-7.9086
1214.000000000,-7.9061
1215.000000000,-7.9035
1216.000000000,-7.9010
1217.000000000,-7.8984
1218.000000000,-7.8959
1219.000000000,-7.8933
1220.000000000,-7.8908
1221.000000000,-7.8882
1222.000000000,-7.8857
1223.000000000,-7.8831
1224.000000000,-7.8806
1225.000000000,-7.8787
1226.000000000,-7.8762
1227.000000000,-7.8737
1228.000000000,-7.8711
1229.000000000,-7.8687
1230.000000000,-7.8662
1231.000000000,-7.8648
1232.000000000,-7.8630
1233.000000000,-7.8605
1234.000000000,-7.8606
1235.000000000,-7.8650
1236.000000000,-7.8639
1237.000000000,-7.8613
1238.000000000,-7.8588
1239.000000000,-7.8563
1240.000000000,-7.8538
1241.000000000,-7.8513
1242.000000000,-7.8488
1243.000000000,-7.8463
1244.000000000,-7.8438
1245.000000000,-7.8414
1246.000000000,-7.8392
1247.000000000,-7.8367
1248.000000000,-7.8350
1249.000000000,-7.8467
1250.000000000,-7.8473
1251.000000000,-7.8451
1252.000000000,-7.8426
1253.000000000,-7.8401
1254.000000000,-7.8376
1255.000000000,-7.8351
1256.000000000,-7.8326
1257.000000000,-7.8301
1258.000000000,-7.8276
1259.000000000,-7.8252
1260.000000000,-7.8228
1261.000000000,-7.8204
1262.000000000,-7.8179
1263.000000000,-7.8154
1264.000000000,-7.8130
1265.000000000,-7.8105
1266.000000000,-7.8081
1267.000000000,-7.8087
1268.000000000,-7.8063
1269.000000000,-7.8038
1270.000000000,-7.8014
1271.000000000,-7.7990
1272.000000000,-7.7965
1273.000000000,-7.7971
1274.000000000,-7.8184
1275.000000000,-7.8168
1276.000000000,-7.8146
1277.000000000,-7.8121
1278.000000000,-7.8096
1279.000000000,-7.8072
1280.000000000,-7.8047
1281.000000000,-7.8022
1282.000000000,-7.7998
1283.000000000,-7.7973
1284.000000000,-7.7949
1285.000000000,-7.7924
1286.000000000,-7.7900
1287.000000000,-7.7876
1288.000000000,-7.7852
1289.000000000,-7.7827
1290.000000000,-7.7803
1291.000000000,-7.7779
1292.000000000,-7.7755
1293.000000000,-7.7730
1294.000000000,-7.7706
1295.000000000,-7.7682
1296.000000000,-7.7658
1297.000000000,-7.7634
1298.000000000,-7.7610
1299.000000000,-7.7586
1300.000000000,-7.7562
1301.000000000,-7.7538
1302.000000000,-7.7515
1303.000000000,-7.7492
1304.000000000,-7.7493
1305.000000000,-7.7471
1306.000000000,-7.7447
1307.000000000,-7.7425
1308.000000000,-7.7401
1309.000000000,-7.7377
1310.000000000,-7.7354
1311.000000000,-7.7330
1312.000000000,-7.7307
1313.000000000,-7.7283
1314.000000000,-7.7260
1315.000000000,-7.7236
1316.000000000,-7.7213
1317.000000000,-7.7190
1318.000000000,-7.7166
1319.000000000,-7.7143
1320.000000000,-7.7120
1321.000000000,-7.7184
1322.000000000,-7.7236
1323.000000000,-7.7241
1324.000000000,-7.7223
1325.000000000,-7.7253
1326.000000000,-7.7246
1327.000000000,-7.7228
1328.000000000,-7.7388
1329.000000000,-7.7387
1330.000000000,-7.7399
1331.000000000,-7.7418
1332.000000000,-7.7394
1333.000000000,-7.7376
1334.000000000,-7.7352
1335.000000000,-7.7328
1336.000000000,-7.7307
1337.000000000,-7.7297
1338.000000000,-7.7279
1339.000000000,-7.7268
1340.000000000,-7.7251
1341.000000000,-7.7235
1342.000000000,-7.7237
1343.000000000,-7.7214
1344.000000000,-7.7190
1345.000000000,-7.7167
1346.000000000,-7.7143
1347.000000000,-7.7120
1348.000000000,-7.7096
1349.000000000,-7.7073
1350.000000000,-7.7059
1351.000000000,-7.7035
1352.000000000,-7.7036
1353.000000000,-7.7014
1354.000000000,-7.7002
1355.000000000,-7.6978
1356.000000000,-7.6955
1357.000000000,-7.6932
1358.000000000,-7.6908
1359.000000000,-7.6885
1360.000000000,-7.6862
1361.000000000,-7.6839
1362.000000000,-7.6816
1363.000000000,-7.6793
1364.000000000,-7.6885
1365.000000000,-7.7125
1366.000000000,-7.7130
1367.000000000,-7.7107
1368.000000000,-7.7083
1369.000000000,-7.7059
1370.000000000,-7.7036
1371.000000000,-7.7012
1372.000000000,-7.6988
1373.000000000,-7.6965
1374.000000000,-7.6941
1375.000000000,-7.6918
1376.000000000,-7.6894
1377.000000000,-7.6872
1378.000000000,-7.6848
1379.000000000,-7.6825
1380.000000000,-7.6802
1381.000000000,-7.6778
1382.000000000,-7.6755
1383.000000000,-7.6732
1384.000000000,-7.6709
1385.000000000,-7.6686
1386.000000000,-7.6663
1387.000000000,-7.6639
1388.000000000,-7.6616
1389.000000000,-7.6594
1390.000000000,-7.6571
1391.000000000,-7.6548
1392.000000000,-7.6525
1393.000000000,-7.6502
1394.000000000,-7.6480
1395.000000000,-7.6457
1396.000000000,-7.6434
1397.000000000,-7.6411
1398.000000000,-7.6389
1399.000000000,-7.6366
1400.000000000,-7.6344
1401.000000000,-7.6321
1402.000000000,-7.6299
1403.000000000,-7.6276
1404.000000000,-7.6304
1405.000000000,-7.6283
1406.000000000,-7.6262
1407.000000000,-7.6246
1408.000000000,-7.6223
1409.000000000,-7.6201
1410.000000000,-7.6254
1411.000000000,-7.6234
1412.000000000,-7.6212
1413.000000000,-7.6189
1414.000000000,-7.6167
1415.000000000,-7.6145
1416.000000000,-7.6122
1417.000000000,-7.6100
1418.000000000,-7.6078
1419.000000000,-7.6056
1420.000000000,-7.6033
1421.000000000,-7.6011
1422.000000000,-7.5989
1423.000000000,-7.5967
1424.000000000,-7.5945
1425.000000000,-7.5923
1426.000000000,-7.5908
1427.000000000,-7.5886
1428.000000000,-7.5864
1429.000000000,-7.5842
1430.000000000,-7.5820
1431.000000000,-7.5799
1432.000000000,-7.5777
1433.000000000,-7.5784
1434.000000000,-7.5811
1435.000000000,-7.5954
1436.000000000,-7.5948
1437.000000000,-7.5926
1438.000000000,-7.5904
1439.000000000,-7.5882
1440.000000000,-7.5860
1441.000000000,-7.5838
1442.000000000,-7.5816
1443.000000000,-7.5798
1444.000000000,-7.5776
1445.000000000,-7.5754
1446.000000000,-7.5733
1447.000000000,-7.5711
1448.000000000,-7.5689
1449.000000000,-7.5668
1450.000000000,-7.5646
1451.000000000,-7.5624
1452.000000000,-7.5606
1453.000000000,-7.5585
1454.000000000,-7.5570
1455.000000000,-7.5548
1456.000000000,-7.5527
1457.000000000,-7.5505
1458.000000000,-7.5484
1459.000000000,-7.5462
1460.000000000,-7.5443
1461.000000000,-7.5422
1462.000000000,-7.5400
1463.000000000,-7.5383
1464.000000000,-7.5362
1465.000000000,-7.5341
1466.000000000,-7.5319
1467.000000000,-7.5298
1468.000000000,-7.5277
1469.000000000,-7.5256
1470.000000000,-7.5235
1471.000000000,-7.5214
1472.000000000,-7.5193
1473.000000000,-7.5172
1474.000000000,-7.5151
1475.000000000,-7.5136
1476.000000000,-7.5128
1477.000000000,-7.5134
1478.000000000,-7.5113
1479.000000000,-7.5127
1480.000000000,-7.5106
1481.000000000,-7.5085
1482.000000000,-7.5064
1483.000000000,-7.5043
1484.000000000,-7.5022
1485.000000000,-7.5002
1486.000000000,-7.4981
1487.000000000,-7.4960
1488.000000000,-7.4940
1489.000000000,-7.4921
1490.000000000,-7.4900
1491.000000000,-7.4880
1492.000000000,-7.4859
1493.000000000,-7.4839
1494.000000000,-7.4818
1495.000000000,-7.4798
1496.000000000,-7.4777
1497.000000000,-7.4758
1498.000000000,-7.4738
1499.000000000,-7.4717
1500.000000000,-7.4697
1501.000000000,-7.4677
1502.000000000,-7.4656
1503.000000000,-7.4636
1504.000000000,-7.4616
1505.000000000,-7.4596
1506.000000000,-7.4688
1507.000000000,-7.4668
1508.000000000,-7.4647
1509.000000000,-7.4629
1510.000000000,-7.4609
1511.000000000,-7.4589
1512.000000000,-7.4583
1513.000000000,-7.4563
1514.000000000,-7.4543
1515.000000000,-7.4523
1516.000000000,-7.4503
1517.000000000,-7.4483
1518.000000000,-7.4463
1519.000000000,-7.4443
1520.000000000,-7.4423
1521.000000000,-7.4403
1522.000000000,-7.4383
1523.000000000,-7.4363
1524.000000000,-7.4343
1525.000000000,-7.4331
1526.000000000,-7.4311
1527.000000000,-7.4292
1528.000000000,-7.4272
1529.000000000,-7.4252
1530.000000000,-7.4233
1531.000000000,-7.4215
1532.000000000,-7.4195
1533.000000000,-7.4176
1534.000000000,-7.4156
1535.000000000,-7.4137
1536.000000000,-7.4117
1537.000000000,-7.4098
1538.000000000,-7.4078
1539.000000000,-7.4059
1540.000000000,-7.4040
1541.000000000,-7.4020
1542.000000000,-7.4001
1543.000000000,-7.3982
1544.000000000,-7.3964
1545.000000000,-7.3945
1546.000000000,-7.3925
1547.000000000,-7.3906
1548.000000000,-7.3887
1549.000000000,-7.3918
1550.000000000,-7.3898
1551.000000000,-7.3879
1552.000000000,-7.3860
1553.000000000,-7.3936
1554.000000000,-7.3916
1555.000000000,-7.3897
1556.000000000,-7.3878
1557.000000000,-7.3859
1558.000000000,-7.3840
1559.000000000,-7.3820
1560.000000000,-7.3801
1561.000000000,-7.3782
1562.000000000,-7.3794
1563.000000000,-7.3783
1564.000000000,-7.3774
1565.000000000,-7.3797
1566.000000000,-7.3778
1567.000000000,-7.3762
1568.000000000,-7.3757
1569.000000000,-7.3738
1570.000000000,-7.3719
1571.000000000,-7.3700
1572.000000000,-7.3681
1573.000000000,-7.3663
1574.000000000,-7.3644
1575.000000000,-7.3625
1576.000000000,-7.3606
1577.000000000,-7.3587
1578.000000000,-7.3568
1579.000000000,-7.3550
1580.000000000,-7.3531
1581.000000000,-7.3512
1582.000000000,-7.3493
1583.000000000,-7.3475
1584.000000000,-7.3456
1585.000000000,-7.3438
1586.000000000,-7.3419
1587.000000000,-7.3400
1588.000000000,-7.3382
1589.000000000,-7.3363
1590.000000000,-7.3345
1591.000000000,-7.3327
1592.000000000,-7.3347
1593.000000000,-7.3329
1594.000000000,-7.3311
1595.000000000,-7.3292
1596.000000000,-7.3274
1597.000000000,-7.3255
1598.000000000,-7.3238
1599.000000000,-7.3220
1600.000000000,-7.3202
1601.000000000,-7.3260
1602.000000000,-7.3247
1603.000000000,-7.3292
1604.000000000,-7.3274
1605.000000000,-7.3258
1606.000000000,-7.3240
1607.000000000,-7.3221
1608.000000000,-7.3203
1609.000000000,-7.3185
1610.000000000,-7.3243
1611.000000000,-7.3226
1612.000000000,-7.3460
1613.000000000,-7.3470
1614.000000000,-7.3457
1615.000000000,-7.3456
1616.000000000,-7.3480
1617.000000000,-7.3467
1618.000000000,-7.3448
1619.000000000,-7.3429
1620.000000000,-7.3410
1621.000000000,-7.3391
1622.000000000,-7.3373
1623.000000000,-7.3354
1624.000000000,-7.3335
1625.000000000,-7.3316
1626.000000000,-7.3298
1627.000000000,-7.3279
1628.000000000,-7.3261
1629.000000000,-7.3242
1630.000000000,-7.3223
1631.000000000,-7.3205
1632.000000000,-7.3186
1633.000000000,-7.3168
1634.000000000,-7.3149
1635.000000000,-7.3131
1636.000000000,-7.3113
1637.000000000,-7.3095
1638.000000000,-7.3077
1639.000000000,-7.3080
1640.000000000,-7.3066
1641.000000000,-7.3047
1642.000000000,-7.3029
1643.000000000,-7.3011
1644.000000000,-7.2993
1645.000000000,-7.2974
1646.000000000,-7.2956
1647.000000000,-7.2941
1648.000000000,-7.2926
1649.000000000,-7.2937
1650.000000000,-7.2956
1651.000000000,-7.2937
1652.000000000,-7.2919
1653.000000000,-7.2901
1654.000000000,-7.2883
1655.000000000,-7.2865
1656.000000000,-7.2853
1657.000000000,-7.2849
1658.000000000,-7.2852
1659.000000000,-7.2843
1660.000000000,-7.2830
1661.000000000,-7.2815
1662.000000000,-7.2797
1663.000000000,-7.2779
1664.000000000,-7.2761
1665.000000000,-7.2744
1666.000000000,-7.2799
1667.000000000,-7.2782
1668.000000000,-7.2764
1669.000000000,-7.2746
1670.000000000,-7.2728
1671.000000000,-7.2710
1672.000000000,-7.2692
1673.000000000,-7.2683
1674.000000000,-7.2669
1675.000000000,-7.2664
1676.000000000,-7.2660
1677.000000000,-7.2642
1678.000000000,-7.2626
1679.000000000,-7.2608
1680.000000000,-7.2590
1681.000000000,-7.2577
1682.000000000,-7.2654
1683.000000000,-7.2636
1684.000000000,-7.2619
1685.000000000,-7.2601
1686.000000000,-7.2583
1687.000000000,-7.2566
1688.000000000,-7.2548
1689.000000000,-7.2537
1690.000000000,-7.2522
1691.000000000,-7.2505
1692.000000000,-7.2487
1693.000000000,-7.2470
1694.000000000,-7.2452
1695.000000000,-7.2434
1696.000000000,-7.2417
1697.000000000,-7.2423
1698.000000000,-7.2433
1699.000000000,-7.2419
1700.000000000,-7.2420
1701.000000000,-7.2402
1702.000000000,-7.2385
1703.000000000,-7.2367
1704.000000000,-7.2350
1705.000000000,-7.2332
1706.000000000,-7.2315
1707.000000000,-7.2297
1708.000000000,-7.2281
1709.000000000,-7.2264
1710.000000000,-7.2247
1711.000000000,-7.2229
1712.000000000,-7.2212
1713.000000000,-7.2195
1714.000000000,-7.2178
1715.000000000,-7.2160
1716.000000000,-7.2143
1717.000000000,-7.2126
1718.000000000,-7.2109
1719.000000000,-7.2092
1720.000000000,-7.2075
1721.000000000,-7.2058
1722.000000000,-7.2040
1723.000000000,-7.2023
1724.000000000,-7.2008
1725.000000000,-7.1991
1726.000000000,-7.1974
1727.000000000,-7.1959
1728.000000000,-7.1942
1729.000000000,-7.2008
1730.000000000,-7.2039
1731.000000000,-7.2189
1732.000000000,-7.2335
1733.000000000,-7.2391
1734.000000000,-7.2396
1735.000000000,-7.2386
1736.000000000,-7.2368
1737.000000000,-7.2350
1738.000000000,-7.2381
1739.000000000,-7.2371
1740.000000000,-7.2353
1741.000000000,-7.2335
1742.000000000,-7.2317
1743.000000000,-7.2300
1744.000000000,-7.2307
1745.000000000,-7.2291
1746.000000000,-7.2273
1747.000000000,-7.2256
1748.000000000,-7.2238
1749.000000000,-7.2220
1750.000000000,-7.2203
1751.000000000,-7.2185
1752.000000000,-7.2168
1753.000000000,-7.2150
1754.000000000,-7.2133
1755.000000000,-7.2115
1756.000000000,-7.2098
1757.000000000,-7.2080
1758.000000000,-7.2063
1759.000000000,-7.2046
1760.000000000,-7.2028
1761.000000000,-7.2011
1762.000000000,-7.1994
1763.000000000,-7.1976
1764.000000000,-7.1959
1765.000000000,-7.1942
1766.000000000,-7.1925
1767.000000000,-7.1908
1768.000000000,-7.1891
1769.000000000,-7.1874
1770.000000000,-7.1857
1771.000000000,-7.1840
1772.000000000,-7.1823
1773.000000000,-7.1806
1774.000000000,-7.1790
1775.000000000,-7.1773
1776.000000000,-7.1756
1777.000000000,-7.1746
1778.000000000,-7.1729
1779.000000000,-7.1715
1780.000000000,-7.1698
1781.000000000,-7.1681
1782.000000000,-7.1664
1783.000000000,-7.1647
1784.000000000,-7.1631
1785.000000000,-7.1614
1786.000000000,-7.1597
1787.000000000,-7.1581
1788.000000000,-7.1564
1789.000000000,-7.1547
1790.000000000,-7.1531
1791.000000000,-7.1514
1792.000000000,-7.1498
1793.000000000,-7.1481
1794.000000000,-7.1465
1795.000000000,-7.1448
1796.000000000,-7.1432
1797.000000000,-7.1415
1798.000000000,-7.1399
1799.000000000,-7.1382
1800.000000000,-7.1366
1801.000000000,-7.1372
1802.000000000,-7.1437
1803.000000000,-7.1443
1804.000000000,-7.1426
1805.000000000,-7.1410
1806.000000000,-7.1393
1807.000000000,-7.1377
1808.000000000,-7.1360
1809.000000000,-7.1344
1810.000000000,-7.1328
1811.000000000,-7.1315
1812.000000000,-7.1327
1813.000000000,-7.1311
1814.000000000,-7.1300
1815.000000000,-7.1284
1816.000000000,-7.1268
1817.000000000,-7.1252
1818.000000000,-7.1236
1819.000000000,-7.1220
1820.000000000,-7.1204
1821.000000000,-7.1188
1822.000000000,-7.1175
1823.000000000,-7.1160
1824.000000000,-7.1144
1825.000000000,-7.1128
1826.000000000,-7.1112
1827.000000000,-7.1096
1828.000000000,-7.1081
1829.000000000,-7.1065
1830.000000000,-7.1049
1831.000000000,-7.1033
1832.000000000,-7.1017
1833.000000000,-7.1001
1834.000000000,-7.0986
1835.000000000,-7.0970
1836.000000000,-7.0954
1837.000000000,-7.0938
1838.000000000,-7.0922
1839.000000000,-7.0907
1840.000000000,-7.0891
1841.000000000,-7.0875
1842.000000000,-7.0861
1843.000000000,-7.0845
1844.000000000,-7.0830
1845.000000000,-7.0816
1846.000000000,-7.0801
1847.000000000,-7.0785
1848.000000000,-7.0770
1849.000000000,-7.0754
1850.000000000,-7.0739
1851.000000000,-7.0723
1852.000000000,-7.0708
1853.000000000,-7.0692
1854.000000000,-7.0677
1855.000000000,-7.0662
1856.000000000,-7.0646
1857.000000000,-7.0631
1858.000000000,-7.0616
1859.000000000,-7.0600
1860.000000000,-7.0587
1861.000000000,-7.0572
1862.000000000,-7.0556
1863.000000000,-7.0541
1864.000000000,-7.0527
1865.000000000,-7.0512
1866.000000000,-7.0497
1867.000000000,-7.0481
1868.000000000,-7.0466
1869.000000000,-7.0451
1870.000000000,-7.0442
1871.000000000,-7.0429
1872.000000000,-7.0414
1873.000000000,-7.0399
1874.000000000,-7.0384
1875.000000000,-7.0369
1876.000000000,-7.0362
1877.000000000,-7.0370
1878.000000000,-7.0449
1879.000000000,-7.0441
1880.000000000,-7.0426
1881.000000000,-7.0413
1882.000000000,-7.0398
1883.000000000,-7.0383
1884.000000000,-7.0368
1885.000000000,-7.0353
1886.000000000,-7.0343
1887.000000000,-7.0328
1888.000000000,-7.0313
1889.000000000,-7.0298
1890.000000000,-7.0283
1891.000000000,-7.0269
1892.000000000,-7.0254
1893.000000000,-7.0239
1894.000000000,-7.0224
1895.000000000,-7.0209
1896.000000000,-7.0195
1897.000000000,-7.0180
1898.000000000,-7.0165
1899.000000000,-7.0150
1900.000000000,-7.0136
1901.000000000,-7.0121
1902.000000000,-7.0107
1903.000000000,-7.0092
1904.000000000,-7.0077
1905.000000000,-7.0063
1906.000000000,-7.0048
1907.000000000,-7.0034
1908.000000000,-7.0019
1909.000000000,-7.0005
1910.000000000,-6.9990
1911.000000000,-6.9976
1912.000000000,-6.9961
1913.000000000,-6.9952
1914.000000000,-6.9937
1915.000000000,-6.9923
1916.000000000,-6.9909
1917.000000000,-6.9894
1918.000000000,-6.9880
1919.000000000,-6.9866
1920.000000000,-6.9851
1921.000000000,-6.9837
1922.000000000,-6.9823
1923.000000000,-6.9809
1924.000000000,-6.9795
1925.000000000,-6.9781
1926.000000000,-6.9766
1927.000000000,-6.9752
1928.000000000,-6.9738
1929.000000000,-6.9724
1930.000000000,-6.9713
1931.000000000,-6.9699
1932.000000000,-6.9685
1933.000000000,-6.9671
1934.000000000,-6.9657
1935.000000000,-6.9643
1936.000000000,-6.9629
1937.000000000,-6.9615
1938.000000000,-6.9603
1939.000000000,-6.9589
1940.000000000,-6.9575
1941.000000000,-6.9561
1942.000000000,-6.9563
1943.000000000,-6.9549
1944.000000000,-6.9535
1945.000000000,-6.9522
1946.000000000,-6.9508
1947.000000000,-6.9494
1948.000000000,-6.9480
1949.000000000,-6.9471
1950.000000000,-6.9566
1951.000000000,-6.9569
1952.000000000,-6.9555
1953.000000000,-6.9541
1954.000000000,-6.9527
1955.000000000,-6.9513
1956.000000000,-6.9499
1957.000000000,-6.9486
1958.000000000,-6.9472
1959.000000000,-6.9458
1960.000000000,-6.9444
1961.000000000,-6.9431
1962.000000000,-6.9417
1963.000000000,-6.9403
1964.000000000,-6.9390
1965.000000000,-6.9377
1966.000000000,-6.9373
1967.000000000,-6.9463
1968.000000000,-6.9451
1969.000000000,-6.9438
1970.000000000,-6.9424
1971.000000000,-6.9410
1972.000000000,-6.9396
1973.000000000,-6.9383
1974.000000000,-6.9369
1975.000000000,-6.9355
1976.000000000,-6.9342
1977.000000000,-6.9328
1978.000000000,-6.9314
1979.000000000,-6.9301
1980.000000000,-6.9287
1981.000000000,-6.9279
1982.000000000,-6.9266
1983.000000000,-6.9252
1984.000000000,-6.9238
1985.000000000,-6.9225
1986.000000000,-6.9212
1987.000000000,-6.9198
1988.000000000,-6.9185
1989.000000000,-6.9172
1990.000000000,-6.9158
1991.000000000,-6.9145
1992.000000000,-6.9131
1993.000000000,-6.9118
1994.000000000,-6.9105
1995.000000000,-6.9092
1996.000000000,-6.9086
1997.000000000,-6.9073
1998.000000000,-6.9059
1999.000000000,-6.9047
2000.000000000,-6.9034
2001.000000000,-6.9021
2002.000000000,-6.9008
2003.000000000,-6.8995
2004.000000000,-6.8982
2005.000000000,-6.8969
2006.000000000,-6.8956
2007.000000000,-6.8948
2008.000000000,-6.8935
2009.000000000,-6.8922
2010.000000000,-6.8909
2011.000000000,-6.8896
2012.000000000,-6.8894
2013.000000000,-6.8900
2014.000000000,-6.8931
2015.000000000,-6.8965
2016.000000000,-6.8971
2017.000000000,-6.8991
2018.000000000,-6.8977
2019.000000000,-6.8964
2020.000000000,-6.8951
2021.000000000,-6.8938
2022.000000000,-6.8925
2023.000000000,-6.8912
2024.000000000,-6.8899
2025.000000000,-6.8885
2026.000000000,-6.8872
2027.000000000,-6.8859
2028.000000000,-6.8846
2029.000000000,-6.8833
2030.000000000,-6.8820
2031.000000000,-6.8807
2032.000000000,-6.8794
2033.000000000,-6.8781
2034.000000000,-6.8768
2035.000000000,-6.8756
2036.000000000,-6.8743
2037.000000000,-6.8730
2038.000000000,-6.8823
2039.000000000,-6.8813
2040.000000000,-6.8800
2041.000000000,-6.8787
2042.000000000,-6.8774
2043.000000000,-6.8761
2044.000000000,-6.8748
2045.000000000,-6.8735
2046.000000000,-6.8722
2047.000000000,-6.8709
2048.000000000,-6.8697
2049.000000000,-6.8724
2050.000000000,-6.8740
2051.000000000,-6.8764
2052.000000000,-6.8760
2053.000000000,-6.8747
2054.000000000,-6.8734
2055.000000000,-6.8721
2056.000000000,-6.8708
2057.000000000,-6.8695
2058.000000000,-6.8691
2059.000000000,-6.8695
2060.000000000,-6.8682
2061.000000000,-6.8669
2062.000000000,-6.8656
2063.000000000,-6.8643
2064.000000000,-6.8630
2065.000000000,-6.8617
2066.000000000,-6.8604
2067.000000000,-6.8592
2068.000000000,-6.8579
2069.000000000,-6.8566
