time,EAST,NORTH,WEST,PATH
1.000000000000,5572.9,2414.0,-15212.,25589.
2.000000000000,5571.3,2413.4,-15258.,25587.
3.000000000000,5568.8,2412.3,-15295.,25584.
4.000000000000,5565.6,2410.8,-15322.,25581.
5.000000000000,5561.7,2409.1,-15337.,25577.
6.000000000000,5557.5,2407.1,-15344.,25572.
7.000000000000,5553.1,2405.0,-15345.,25568.
8.000000000000,5548.6,2402.7,-15341.,25563.
9.000000000000,5544.1,2400.3,-15340.,25559.
10.00000000000,5539.7,2397.9,-15340.,25555.
11.00000000000,5535.3,2395.5,-15331.,25552.
12.00000000000,5531.1,2393.0,-15316.,25548.
13.00000000000,5526.9,2390.5,-15301.,25545.
14.00000000000,5522.9,2388.0,-15285.,25542.
15.00000000000,5519.1,2385.6,-15270.,25539.
16.00000000000,5515.4,2383.2,-15255.,25537.
17.00000000000,5511.9,2380.8,-15240.,25535.
18.00000000000,5508.5,2378.5,-15225.,25532.
19.00000000000,5505.3,2376.2,-15210.,25530.
20.00000000000,5502.3,2373.9,-15196.,25529.
21.00000000000,5499.4,2371.7,-15181.,25527.
22.00000000000,5496.6,2369.6,-15167.,25525.
23.00000000000,5493.9,2367.5,-15152.,25524.
24.00000000000,5491.3,2365.5,-15138.,25522.
25.00000000000,5488.9,2363.5,-15124.,25521.
26.00000000000,5486.4,2361.5,-15110.,25520.
27.00000000000,5484.1,2359.7,-15096.,25518.
28.00000000000,5481.9,2357.8,-15082.,25517.
29.00000000000,5479.7,2356.1,-15068.,25516.
30.00000000000,5477.6,2354.4,-15055.,25515.
31.00000000000,5475.6,2352.8,-15041.,25514.
32.00000000000,5473.8,2351.3,-15027.,25513.
33.00000000000,5472.0,2349.8,-15014.,25512.
34.00000000000,5470.2,2348.4,-15001.,25511.
35.00000000000,5468.6,2347.0,-14987.,25510.
36.00000000000,5467.1,2345.8,-14974.,25509.
37.00000000000,5465.6,2344.5,-14961.,25508.
38.00000000000,5464.2,2343.3,-14948.,25507.
39.00000000000,5462.9,2342.2,-14935.,25507.
40.00000000000,5461.7,2341.1,-14923.,25506.
41.00000000000,5460.5,2340.1,-14910.,25505.
42.00000000000,5459.4,2339.1,-14898.,25505.
43.00000000000,5458.4,2338.2,-14886.,25504.
44.00000000000,5457.4,2337.3,-14874.,25504.
45.00000000000,5456.5,2336.5,-14862.,25503.
46.00000000000,5455.6,2335.6,-14850.,25503.
47.00000000000,5454.8,2334.9,-14839.,25502.
48.00000000000,5454.0,2334.1,-14827.,25502.
49.00000000000,5453.3,2333.4,-14816.,25501.
50.00000000000,5452.6,2332.7,-14805.,25501.
51.00000000000,5451.9,2332.1,-14794.,25501.
52.00000000000,5451.3,2331.4,-14783.,25500.
53.00000000000,5450.7,2330.9,-14772.,25500.
54.00000000000,5450.2,2330.3,-14762.,25500.
55.00000000000,5449.7,2329.7,-14751.,25499.
56.00000000000,5449.2,2329.2,-14740.,25499.
57.00000000000,5448.7,2328.7,-14730.,25499.
58.00000000000,5448.2,2328.2,-14720.,25498.
59.00000000000,5447.8,2327.7,-14709.,25498.
60.00000000000,5447.4,2327.3,-14699.,25498.
61.00000000000,5447.0,2326.9,-14689.,25497.
62.00000000000,5446.6,2326.4,-14679.,25497.
63.00000000000,5446.2,2326.0,-14669.,25497.
64.00000000000,5445.8,2325.6,-14659.,25496.
65.00000000000,5445.5,2325.3,-14650.,25496.
66.00000000000,5445.2,2324.9,-14640.,25496.
67.00000000000,5444.8,2324.5,-14631.,25495.
68.00000000000,5444.4,2324.2,-14621.,25495.
69.00000000000,5444.0,2323.9,-14612.,25495.
70.00000000000,5443.6,2323.6,-14603.,25495.
71.00000000000,5443.1,2323.2,-14594.,25494.
72.00000000000,5442.6,2322.9,-14584.,25494.
73.00000000000,5442.1,2322.7,-14575.,25494.
74.00000000000,5441.6,2322.4,-14566.,25493.
75.00000000000,5441.3,2322.1,-14557.,25493.
76.00000000000,5440.9,2321.8,-14548.,25493.
77.00000000000,5440.6,2321.6,-14539.,25493.
78.00000000000,5440.3,2321.3,-14530.,25492.
79.00000000000,5440.0,2321.1,-14521.,25492.
80.00000000000,5439.7,2320.8,-14513.,25492.
81.00000000000,5439.5,2320.6,-14504.,25491.
82.00000000000,5439.2,2320.3,-14496.,25491.
83.00000000000,5439.0,2320.1,-14487.,25491.
84.00000000000,5438.7,2319.9,-14479.,25491.
85.00000000000,5438.5,2319.7,-14470.,25490.
86.00000000000,5438.3,2319.5,-14462.,25490.
87.00000000000,5438.1,2319.2,-14453.,25490.
88.00000000000,5437.9,2319.0,-14445.,25490.
89.00000000000,5437.7,2318.8,-14437.,25489.
90.00000000000,5437.5,2318.6,-14428.,25489.
91.00000000000,5437.3,2318.4,-14420.,25489.
92.00000000000,5437.2,2318.2,-14412.,25489.
93.00000000000,5437.0,2318.1,-14405.,25489.
94.00000000000,5436.8,2317.9,-14398.,25488.
95.00000000000,5436.6,2317.7,-14390.,25488.
96.00000000000,5436.5,2317.5,-14381.,25488.
97.00000000000,5436.3,2317.3,-14373.,25488.
98.00000000000,5436.1,2317.1,-14365.,25487.
99.00000000000,5436.0,2317.0,-14357.,25487.
100.0000000000,5435.8,2316.8,-14349.,25487.
101.0000000000,5435.6,2316.6,-14342.,25487.
102.0000000000,5435.5,2316.4,-14334.,25486.
103.0000000000,5435.3,2316.3,-14326.,25486.
104.0000000000,5435.2,2316.1,-14318.,25486.
105.0000000000,5435.0,2315.9,-14311.,25486.
106.0000000000,5434.9,2315.8,-14303.,25486.
107.0000000000,5434.7,2315.6,-14296.,25485.
108.0000000000,5434.6,2315.5,-14289.,25485.
109.0000000000,5434.4,2315.3,-14282.,25485.
110.0000000000,5434.3,2315.1,-14274.,25485.
111.0000000000,5434.1,2315.0,-14266.,25485.
112.0000000000,5434.0,2314.8,-14259.,25484.
113.0000000000,5433.8,2314.7,-14251.,25484.
114.0000000000,5433.7,2314.5,-14244.,25484.
115.0000000000,5433.5,2314.4,-14237.,25484.
116.0000000000,5433.4,2314.2,-14229.,25484.
117.0000000000,5433.3,2314.1,-14222.,25483.
118.0000000000,5433.1,2313.9,-14217.,25483.
119.0000000000,5433.0,2313.8,-14215.,25483.
120.0000000000,5432.8,2313.6,-14209.,25483.
121.0000000000,5432.7,2313.5,-14201.,25483.
122.0000000000,5432.6,2313.3,-14194.,25482.
123.0000000000,5432.4,2313.2,-14187.,25482.
124.0000000000,5432.3,2313.0,-14179.,25482.
125.0000000000,5432.2,2312.9,-14171.,25482.
126.0000000000,5432.0,2312.8,-14164.,25482.
127.0000000000,5431.9,2312.6,-14157.,25482.
128.0000000000,5431.8,2312.5,-14150.,25481.
129.0000000000,5431.6,2312.3,-14143.,25481.
130.0000000000,5431.5,2312.2,-14136.,25481.
131.0000000000,5431.4,2312.1,-14130.,25481.
132.0000000000,5431.2,2311.9,-14124.,25481.
133.0000000000,5431.1,2311.8,-14117.,25480.
134.0000000000,5431.0,2311.7,-14110.,25480.
135.0000000000,5430.8,2311.5,-14104.,25480.
136.0000000000,5430.7,2311.4,-14097.,25480.
137.0000000000,5430.6,2311.2,-14090.,25480.
138.0000000000,5430.5,2311.1,-14083.,25480.
139.0000000000,5430.3,2311.0,-14076.,25479.
140.0000000000,5430.2,2310.8,-14069.,25479.
141.0000000000,5430.1,2310.7,-14063.,25479.
142.0000000000,5430.0,2310.6,-14056.,25479.
143.0000000000,5429.8,2310.4,-14049.,25479.
144.0000000000,5429.7,2310.3,-14045.,25479.
145.0000000000,5429.6,2310.2,-14039.,25478.
146.0000000000,5429.5,2310.1,-14036.,25478.
147.0000000000,5429.4,2309.9,-14031.,25478.
148.0000000000,5429.2,2309.8,-14024.,25478.
149.0000000000,5429.1,2309.7,-14017.,25478.
150.0000000000,5429.0,2309.5,-14010.,25478.
151.0000000000,5428.9,2309.4,-14003.,25477.
152.0000000000,5428.8,2309.3,-13996.,25477.
153.0000000000,5428.7,2309.2,-13989.,25477.
154.0000000000,5428.5,2309.0,-13983.,25477.
155.0000000000,5428.4,2308.9,-13976.,25477.
156.0000000000,5428.3,2308.8,-13970.,25477.
157.0000000000,5428.2,2308.7,-13963.,25476.
158.0000000000,5428.1,2308.6,-13957.,25476.
159.0000000000,5428.0,2308.4,-13951.,25476.
160.0000000000,5427.9,2308.3,-13945.,25476.
161.0000000000,5427.7,2308.2,-13938.,25476.
162.0000000000,5427.6,2308.1,-13932.,25476.
163.0000000000,5427.5,2308.0,-13925.,25476.
164.0000000000,5427.4,2307.8,-13919.,25475.
165.0000000000,5427.3,2307.7,-13913.,25475.
166.0000000000,5427.2,2307.6,-13910.,25475.
167.0000000000,5427.1,2307.5,-13906.,25475.
168.0000000000,5427.0,2307.4,-13900.,25475.
169.0000000000,5426.9,2307.3,-13893.,25475.
170.0000000000,5426.8,2307.2,-13886.,25474.
171.0000000000,5426.7,2307.0,-13880.,25474.
172.0000000000,5426.6,2306.9,-13873.,25474.
173.0000000000,5426.5,2306.8,-13867.,25474.
174.0000000000,5426.4,2306.7,-13860.,25474.
175.0000000000,5426.3,2306.6,-13854.,25474.
176.0000000000,5426.2,2306.5,-13848.,25474.
177.0000000000,5426.1,2306.4,-13841.,25474.
178.0000000000,5426.0,2306.3,-13835.,25473.
179.0000000000,5425.9,2306.2,-13829.,25473.
180.0000000000,5425.8,2306.1,-13823.,25473.
181.0000000000,5425.7,2306.0,-13817.,25473.
182.0000000000,5425.6,2305.9,-13811.,25473.
183.0000000000,5425.5,2305.8,-13805.,25473.
184.0000000000,5425.4,2305.7,-13799.,25473.
185.0000000000,5425.3,2305.6,-13793.,25472.
186.0000000000,5425.2,2305.5,-13787.,25472.
187.0000000000,5425.1,2305.4,-13781.,25472.
188.0000000000,5425.1,2305.3,-13774.,25472.
189.0000000000,5425.0,2305.2,-13768.,25472.
190.0000000000,5424.9,2305.1,-13762.,25472.
191.0000000000,5424.8,2305.1,-13756.,25472.
192.0000000000,5424.7,2305.0,-13750.,25472.
193.0000000000,5424.6,2304.9,-13744.,25472.
194.0000000000,5424.6,2304.8,-13738.,25471.
195.0000000000,5424.5,2304.8,-13731.,25471.
196.0000000000,5424.4,2304.7,-13726.,25471.
197.0000000000,5424.3,2304.6,-13721.,25471.
198.0000000000,5424.3,2304.6,-13717.,25471.
199.0000000000,5424.2,2304.5,-13712.,25471.
200.0000000000,5424.1,2304.4,-13707.,25471.
201.0000000000,5424.1,2304.4,-13700.,25471.
202.0000000000,5424.0,2304.3,-13694.,25471.
203.0000000000,5423.9,2304.3,-13688.,25470.
204.0000000000,5423.9,2304.2,-13682.,25470.
205.0000000000,5423.8,2304.2,-13676.,25470.
206.0000000000,5423.7,2304.1,-13670.,25470.
207.0000000000,5423.7,2304.1,-13664.,25470.
208.0000000000,5423.6,2304.0,-13658.,25470.
209.0000000000,5423.6,2304.0,-13652.,25470.
210.0000000000,5423.5,2303.9,-13646.,25470.
211.0000000000,5423.5,2303.9,-13640.,25470.
212.0000000000,5423.4,2303.8,-13634.,25470.
213.0000000000,5423.4,2303.8,-13629.,25469.
214.0000000000,5423.3,2303.8,-13623.,25469.
215.0000000000,5423.3,2303.7,-13617.,25469.
216.0000000000,5423.2,2303.7,-13611.,25469.
217.0000000000,5423.2,2303.7,-13605.,25469.
218.0000000000,5423.1,2303.6,-13599.,25469.
219.0000000000,5423.1,2303.6,-13593.,25469.
220.0000000000,5423.0,2303.6,-13587.,25469.
221.0000000000,5423.0,2303.5,-13581.,25469.
222.0000000000,5423.0,2303.5,-13575.,25469.
223.0000000000,5422.9,2303.5,-13569.,25469.
224.0000000000,5422.9,2303.4,-13563.,25469.
225.0000000000,5422.9,2303.4,-13558.,25469.
226.0000000000,5422.8,2303.4,-13552.,25468.
227.0000000000,5422.8,2303.4,-13546.,25468.
228.0000000000,5422.8,2303.3,-13540.,25468.
229.0000000000,5422.7,2303.3,-13534.,25468.
230.0000000000,5422.7,2303.3,-13528.,25468.
231.0000000000,5422.7,2303.3,-13522.,25468.
232.0000000000,5422.6,2303.3,-13516.,25468.
233.0000000000,5422.6,2303.2,-13511.,25468.
234.0000000000,5422.6,2303.2,-13505.,25468.
235.0000000000,5422.6,2303.2,-13499.,25468.
236.0000000000,5422.6,2303.2,-13495.,25468.
237.0000000000,5422.5,2303.2,-13490.,25468.
238.0000000000,5422.5,2303.2,-13484.,25468.
239.0000000000,5422.5,2303.2,-13480.,25468.
240.0000000000,5422.5,2303.2,-13477.,25468.
241.0000000000,5422.5,2303.1,-13472.,25468.
242.0000000000,5422.4,2303.1,-13466.,25467.
243.0000000000,5422.4,2303.1,-13460.,25467.
244.0000000000,5422.4,2303.1,-13454.,25467.
245.0000000000,5422.4,2303.1,-13449.,25467.
246.0000000000,5422.3,2303.1,-13443.,25467.
247.0000000000,5422.2,2303.1,-13438.,25467.
248.0000000000,5422.1,2303.1,-13433.,25467.
249.0000000000,5422.0,2303.1,-13428.,25467.
250.0000000000,5422.0,2303.1,-13422.,25467.
251.0000000000,5421.9,2303.1,-13416.,25467.
252.0000000000,5421.9,2303.1,-13411.,25467.
253.0000000000,5421.9,2303.1,-13405.,25467.
254.0000000000,5421.9,2303.1,-13400.,25467.
255.0000000000,5421.9,2303.1,-13394.,25467.
256.0000000000,5421.9,2303.1,-13389.,25467.
257.0000000000,5421.9,2303.1,-13383.,25467.
258.0000000000,5421.9,2303.1,-13377.,25467.
259.0000000000,5421.8,2303.1,-13371.,25467.
260.0000000000,5421.8,2303.1,-13365.,25467.
261.0000000000,5421.8,2303.1,-13360.,25467.
262.0000000000,5421.8,2303.1,-13355.,25467.
263.0000000000,5421.9,2303.1,-13353.,25467.
264.0000000000,5421.9,2303.1,-13352.,25467.
265.0000000000,5421.9,2303.1,-13348.,25467.
266.0000000000,5421.9,2303.1,-13343.,25467.
267.0000000000,5421.9,2303.1,-13337.,25467.
268.0000000000,5421.9,2303.1,-13331.,25467.
269.0000000000,5421.9,2303.2,-13325.,25467.
270.0000000000,5421.9,2303.2,-13320.,25467.
271.0000000000,5421.9,2303.2,-13314.,25466.
272.0000000000,5422.0,2303.2,-13309.,25466.
273.0000000000,5422.0,2303.2,-13303.,25466.
274.0000000000,5422.0,2303.2,-13297.,25466.
275.0000000000,5422.0,2303.2,-13292.,25466.
276.0000000000,5422.0,2303.2,-13286.,25466.
277.0000000000,5422.0,2303.2,-13281.,25466.
278.0000000000,5422.1,2303.2,-13275.,25466.
279.0000000000,5422.1,2303.2,-13270.,25466.
280.0000000000,5422.1,2303.2,-13264.,25466.
281.0000000000,5422.1,2303.3,-13258.,25466.
282.0000000000,5422.2,2303.3,-13253.,25466.
283.0000000000,5422.2,2303.3,-13247.,25466.
284.0000000000,5422.2,2303.3,-13242.,25466.
285.0000000000,5422.2,2303.3,-13236.,25466.
286.0000000000,5422.3,2303.3,-13231.,25466.
287.0000000000,5422.3,2303.3,-13226.,25467.
288.0000000000,5422.3,2303.3,-13221.,25467.
289.0000000000,5422.4,2303.3,-13219.,25467.
290.0000000000,5422.4,2303.3,-13215.,25467.
291.0000000000,5422.4,2303.4,-13210.,25467.
292.0000000000,5422.4,2303.4,-13204.,25467.
293.0000000000,5422.5,2303.4,-13199.,25467.
294.0000000000,5422.5,2303.4,-13193.,25467.
295.0000000000,5422.5,2303.4,-13188.,25467.
296.0000000000,5422.6,2303.4,-13182.,25467.
297.0000000000,5422.6,2303.4,-13177.,25467.
298.0000000000,5422.6,2303.4,-13171.,25467.
299.0000000000,5422.7,2303.4,-13166.,25467.
300.0000000000,5422.7,2303.5,-13161.,25467.
301.0000000000,5422.7,2303.5,-13155.,25467.
302.0000000000,5422.8,2303.5,-13150.,25467.
303.0000000000,5422.8,2303.5,-13145.,25467.
304.0000000000,5422.8,2303.5,-13139.,25467.
305.0000000000,5422.9,2303.5,-13134.,25467.
306.0000000000,5422.9,2303.5,-13128.,25467.
307.0000000000,5423.0,2303.5,-13123.,25467.
308.0000000000,5423.0,2303.5,-13118.,25467.
309.0000000000,5423.0,2303.6,-13113.,25467.
310.0000000000,5423.1,2303.6,-13107.,25467.
311.0000000000,5423.1,2303.6,-13102.,25467.
312.0000000000,5423.1,2303.6,-13097.,25467.
313.0000000000,5423.2,2303.6,-13092.,25467.
314.0000000000,5423.2,2303.6,-13086.,25467.
315.0000000000,5423.3,2303.6,-13081.,25467.
316.0000000000,5423.3,2303.6,-13075.,25467.
317.0000000000,5423.3,2303.7,-13070.,25467.
318.0000000000,5423.4,2303.7,-13064.,25467.
319.0000000000,5423.4,2303.7,-13059.,25467.
320.0000000000,5423.5,2303.7,-13054.,25467.
321.0000000000,5423.5,2303.7,-13048.,25467.
322.0000000000,5423.5,2303.7,-13043.,25468.
323.0000000000,5423.6,2303.7,-13037.,25468.
324.0000000000,5423.6,2303.7,-13032.,25468.
325.0000000000,5423.7,2303.8,-13027.,25468.
326.0000000000,5423.7,2303.8,-13021.,25468.
327.0000000000,5423.7,2303.8,-13016.,25468.
328.0000000000,5423.8,2303.8,-13011.,25468.
329.0000000000,5423.8,2303.8,-13007.,25468.
330.0000000000,5423.9,2303.8,-13002.,25468.
331.0000000000,5423.9,2303.8,-12997.,25468.
332.0000000000,5424.0,2303.8,-12992.,25468.
333.0000000000,5424.0,2303.9,-12986.,25468.
334.0000000000,5424.1,2303.9,-12981.,25468.
335.0000000000,5424.1,2303.9,-12976.,25468.
336.0000000000,5424.1,2303.9,-12970.,25468.
337.0000000000,5424.2,2303.9,-12965.,25468.
338.0000000000,5424.2,2303.9,-12960.,25468.
339.0000000000,5424.3,2303.9,-12955.,25468.
340.0000000000,5424.3,2304.0,-12950.,25468.
341.0000000000,5424.4,2304.0,-12945.,25468.
342.0000000000,5424.4,2304.0,-12939.,25468.
343.0000000000,5424.5,2304.0,-12934.,25469.
344.0000000000,5424.5,2304.0,-12929.,25469.
345.0000000000,5424.6,2304.0,-12924.,25469.
346.0000000000,5424.6,2304.0,-12919.,25469.
347.0000000000,5424.7,2304.0,-12913.,25469.
348.0000000000,5424.7,2304.1,-12908.,25469.
349.0000000000,5424.8,2304.1,-12903.,25469.
350.0000000000,5424.8,2304.1,-12898.,25469.
351.0000000000,5424.9,2304.1,-12893.,25469.
352.0000000000,5424.9,2304.1,-12888.,25469.
353.0000000000,5425.0,2304.1,-12882.,25469.
354.0000000000,5425.0,2304.1,-12877.,25469.
355.0000000000,5425.0,2304.1,-12873.,25469.
356.0000000000,5425.1,2304.2,-12868.,25469.
357.0000000000,5425.1,2304.2,-12863.,25469.
358.0000000000,5425.2,2304.2,-12858.,25469.
359.0000000000,5425.2,2304.2,-12853.,25469.
360.0000000000,5425.2,2304.2,-12848.,25469.
361.0000000000,5425.3,2304.2,-12843.,25470.
362.0000000000,5425.3,2304.2,-12838.,25470.
363.0000000000,5425.4,2304.3,-12834.,25470.
364.0000000000,5425.4,2304.3,-12829.,25470.
365.0000000000,5425.5,2304.3,-12823.,25470.
366.0000000000,5425.5,2304.3,-12818.,25470.
367.0000000000,5425.5,2304.3,-12813.,25470.
368.0000000000,5425.6,2304.3,-12808.,25470.
369.0000000000,5425.6,2304.3,-12803.,25470.
370.0000000000,5425.7,2304.4,-12798.,25470.
371.0000000000,5425.7,2304.4,-12793.,25470.
372.0000000000,5425.8,2304.4,-12788.,25470.
373.0000000000,5425.8,2304.4,-12783.,25470.
374.0000000000,5425.9,2304.4,-12778.,25470.
375.0000000000,5425.9,2304.4,-12773.,25470.
376.0000000000,5426.0,2304.4,-12768.,25470.
377.0000000000,5426.0,2304.4,-12763.,25471.
378.0000000000,5426.1,2304.5,-12758.,25471.
379.0000000000,5426.1,2304.5,-12753.,25471.
380.0000000000,5426.2,2304.5,-12747.,25471.
381.0000000000,5426.2,2304.5,-12742.,25471.
382.0000000000,5426.3,2304.5,-12737.,25471.
383.0000000000,5426.3,2304.5,-12732.,25471.
384.0000000000,5426.4,2304.5,-12727.,25471.
385.0000000000,5426.4,2304.6,-12722.,25471.
386.0000000000,5426.5,2304.6,-12717.,25471.
387.0000000000,5426.5,2304.6,-12712.,25471.
388.0000000000,5426.6,2304.6,-12707.,25471.
389.0000000000,5426.6,2304.6,-12702.,25471.
390.0000000000,5426.7,2304.6,-12697.,25471.
391.0000000000,5426.7,2304.6,-12692.,25471.
392.0000000000,5426.8,2304.7,-12687.,25472.
393.0000000000,5426.8,2304.7,-12682.,25472.
394.0000000000,5426.9,2304.7,-12677.,25472.
395.0000000000,5426.9,2304.7,-12672.,25472.
396.0000000000,5427.0,2304.7,-12667.,25472.
397.0000000000,5427.0,2304.7,-12662.,25472.
398.0000000000,5427.1,2304.7,-12657.,25472.
399.0000000000,5427.1,2304.7,-12652.,25472.
400.0000000000,5427.2,2304.8,-12647.,25472.
401.0000000000,5427.2,2304.8,-12642.,25472.
402.0000000000,5427.3,2304.8,-12638.,25472.
403.0000000000,5427.3,2304.8,-12633.,25472.
404.0000000000,5427.4,2304.8,-12628.,25472.
405.0000000000,5427.4,2304.8,-12623.,25473.
406.0000000000,5427.5,2304.8,-12618.,25473.
407.0000000000,5427.5,2304.9,-12613.,25473.
408.0000000000,5427.6,2304.9,-12608.,25473.
409.0000000000,5427.6,2304.9,-12603.,25473.
410.0000000000,5427.7,2304.9,-12598.,25473.
411.0000000000,5427.7,2304.9,-12593.,25473.
412.0000000000,5427.8,2304.9,-12588.,25473.
413.0000000000,5427.8,2304.9,-12583.,25473.
414.0000000000,5427.9,2305.0,-12578.,25473.
415.0000000000,5427.9,2305.0,-12574.,25473.
416.0000000000,5428.0,2305.0,-12569.,25473.
417.0000000000,5428.0,2305.0,-12564.,25473.
418.0000000000,5428.1,2305.0,-12559.,25474.
419.0000000000,5428.1,2305.0,-12554.,25474.
420.0000000000,5428.2,2305.0,-12549.,25474.
421.0000000000,5428.2,2305.1,-12544.,25474.
422.0000000000,5428.3,2305.1,-12540.,25474.
423.0000000000,5428.3,2305.1,-12535.,25474.
424.0000000000,5428.4,2305.1,-12531.,25474.
425.0000000000,5428.4,2305.1,-12526.,25474.
426.0000000000,5428.5,2305.1,-12521.,25474.
427.0000000000,5428.5,2305.1,-12516.,25474.
428.0000000000,5428.6,2305.2,-12511.,25474.
429.0000000000,5428.6,2305.2,-12507.,25474.
430.0000000000,5428.7,2305.2,-12502.,25475.
431.0000000000,5428.7,2305.2,-12497.,25475.
432.0000000000,5428.8,2305.2,-12492.,25475.
433.0000000000,5428.9,2305.2,-12487.,25475.
434.0000000000,5428.9,2305.2,-12483.,25475.
435.0000000000,5429.0,2305.3,-12478.,25475.
436.0000000000,5429.0,2305.3,-12473.,25475.
437.0000000000,5429.1,2305.3,-12468.,25475.
438.0000000000,5429.1,2305.3,-12464.,25475.
439.0000000000,5429.2,2305.3,-12459.,25475.
440.0000000000,5429.2,2305.3,-12454.,25475.
441.0000000000,5429.3,2305.3,-12449.,25475.
442.0000000000,5429.3,2305.4,-12445.,25476.
443.0000000000,5429.4,2305.4,-12440.,25476.
444.0000000000,5429.4,2305.4,-12435.,25476.
445.0000000000,5429.5,2305.4,-12430.,25476.
446.0000000000,5429.5,2305.4,-12426.,25476.
447.0000000000,5429.6,2305.4,-12421.,25476.
448.0000000000,5429.6,2305.4,-12416.,25476.
449.0000000000,5429.7,2305.5,-12412.,25476.
450.0000000000,5429.7,2305.5,-12407.,25476.
451.0000000000,5429.8,2305.5,-12402.,25476.
452.0000000000,5429.8,2305.5,-12397.,25476.
453.0000000000,5429.9,2305.5,-12393.,25477.
454.0000000000,5429.9,2305.5,-12388.,25477.
455.0000000000,5430.0,2305.5,-12383.,25477.
456.0000000000,5430.0,2305.6,-12379.,25477.
457.0000000000,5430.1,2305.6,-12374.,25477.
458.0000000000,5430.1,2305.6,-12369.,25477.
459.0000000000,5430.2,2305.6,-12365.,25477.
460.0000000000,5430.2,2305.6,-12361.,25477.
461.0000000000,5430.3,2305.6,-12356.,25477.
462.0000000000,5430.3,2305.7,-12351.,25477.
463.0000000000,5430.4,2305.7,-12347.,25477.
464.0000000000,5430.4,2305.7,-12342.,25478.
465.0000000000,5430.5,2305.7,-12337.,25478.
466.0000000000,5430.6,2305.7,-12333.,25478.
467.0000000000,5430.6,2305.7,-12328.,25478.
468.0000000000,5430.7,2305.7,-12324.,25478.
469.0000000000,5430.7,2305.8,-12319.,25478.
470.0000000000,5430.8,2305.8,-12314.,25478.
471.0000000000,5430.8,2305.8,-12310.,25478.
472.0000000000,5430.9,2305.8,-12305.,25478.
473.0000000000,5430.9,2305.8,-12300.,25478.
474.0000000000,5431.0,2305.8,-12296.,25478.
475.0000000000,5431.0,2305.8,-12291.,25479.
476.0000000000,5431.1,2305.9,-12287.,25479.
477.0000000000,5431.1,2305.9,-12282.,25479.
478.0000000000,5431.2,2305.9,-12278.,25479.
479.0000000000,5431.2,2305.9,-12273.,25479.
480.0000000000,5431.3,2305.9,-12268.,25479.
481.0000000000,5431.3,2305.9,-12264.,25479.
482.0000000000,5431.4,2305.9,-12259.,25479.
483.0000000000,5431.4,2306.0,-12255.,25479.
484.0000000000,5431.5,2306.0,-12250.,25479.
485.0000000000,5431.5,2306.0,-12246.,25480.
486.0000000000,5431.6,2306.0,-12241.,25480.
487.0000000000,5431.6,2306.0,-12237.,25480.
488.0000000000,5431.7,2306.0,-12232.,25480.
489.0000000000,5431.8,2306.1,-12227.,25480.
490.0000000000,5431.8,2306.1,-12223.,25480.
491.0000000000,5431.9,2306.1,-12218.,25480.
492.0000000000,5431.9,2306.1,-12214.,25480.
493.0000000000,5432.0,2306.1,-12210.,25480.
494.0000000000,5432.0,2306.1,-12205.,25480.
495.0000000000,5432.1,2306.1,-12201.,25481.
496.0000000000,5432.1,2306.2,-12197.,25481.
497.0000000000,5432.2,2306.2,-12192.,25481.
498.0000000000,5432.2,2306.2,-12188.,25481.
499.0000000000,5432.3,2306.2,-12184.,25481.
500.0000000000,5432.3,2306.2,-12179.,25481.
501.0000000000,5432.4,2306.2,-12175.,25481.
502.0000000000,5432.4,2306.2,-12171.,25481.
503.0000000000,5432.5,2306.3,-12166.,25481.
504.0000000000,5432.5,2306.3,-12162.,25481.
505.0000000000,5432.6,2306.3,-12157.,25482.
506.0000000000,5432.7,2306.3,-12153.,25482.
507.0000000000,5432.7,2306.3,-12148.,25482.
508.0000000000,5432.8,2306.3,-12144.,25482.
509.0000000000,5432.8,2306.4,-12139.,25482.
510.0000000000,5432.9,2306.4,-12135.,25482.
511.0000000000,5432.9,2306.4,-12133.,25482.
512.0000000000,5433.0,2306.4,-12129.,25482.
513.0000000000,5433.0,2306.4,-12125.,25482.
514.0000000000,5433.1,2306.4,-12121.,25482.
515.0000000000,5433.1,2306.4,-12116.,25483.
516.0000000000,5433.2,2306.5,-12112.,25483.
517.0000000000,5433.2,2306.5,-12107.,25483.
518.0000000000,5433.3,2306.5,-12103.,25483.
519.0000000000,5433.3,2306.5,-12099.,25483.
520.0000000000,5433.4,2306.5,-12094.,25483.
521.0000000000,5433.5,2306.5,-12090.,25483.
522.0000000000,5433.5,2306.6,-12085.,25483.
523.0000000000,5433.6,2306.6,-12081.,25483.
524.0000000000,5433.6,2306.6,-12077.,25484.
525.0000000000,5433.7,2306.6,-12072.,25484.
526.0000000000,5433.7,2306.6,-12068.,25484.
527.0000000000,5433.8,2306.6,-12064.,25484.
528.0000000000,5433.8,2306.6,-12059.,25484.
529.0000000000,5433.9,2306.7,-12055.,25484.
530.0000000000,5433.9,2306.7,-12052.,25484.
531.0000000000,5434.0,2306.7,-12048.,25484.
532.0000000000,5434.0,2306.7,-12043.,25484.
533.0000000000,5434.1,2306.7,-12039.,25484.
534.0000000000,5434.1,2306.7,-12035.,25485.
535.0000000000,5434.2,2306.8,-12030.,25485.
536.0000000000,5434.3,2306.8,-12029.,25485.
537.0000000000,5434.3,2306.8,-12028.,25485.
538.0000000000,5434.4,2306.8,-12025.,25485.
539.0000000000,5434.4,2306.8,-12022.,25485.
540.0000000000,5434.5,2306.8,-12018.,25485.
541.0000000000,5434.5,2306.8,-12015.,25485.
542.0000000000,5434.6,2306.9,-12011.,25485.
543.0000000000,5434.6,2306.9,-12007.,25486.
544.0000000000,5434.7,2306.9,-12003.,25486.
545.0000000000,5434.7,2306.9,-11999.,25486.
546.0000000000,5434.8,2306.9,-11994.,25486.
547.0000000000,5434.8,2306.9,-11990.,25486.
548.0000000000,5434.9,2307.0,-11986.,25486.
549.0000000000,5435.0,2307.0,-11982.,25486.
550.0000000000,5435.0,2307.0,-11977.,25486.
551.0000000000,5435.1,2307.0,-11973.,25486.
552.0000000000,5435.1,2307.0,-11969.,25487.
553.0000000000,5435.2,2307.0,-11964.,25487.
554.0000000000,5435.2,2307.0,-11960.,25487.
555.0000000000,5435.3,2307.1,-11956.,25487.
556.0000000000,5435.3,2307.1,-11952.,25487.
557.0000000000,5435.4,2307.1,-11947.,25487.
558.0000000000,5435.4,2307.1,-11943.,25487.
559.0000000000,5435.5,2307.1,-11939.,25487.
560.0000000000,5435.5,2307.1,-11935.,25487.
561.0000000000,5435.6,2307.2,-11931.,25488.
562.0000000000,5435.7,2307.2,-11927.,25488.
563.0000000000,5435.7,2307.2,-11923.,25488.
564.0000000000,5435.8,2307.2,-11919.,25488.
565.0000000000,5435.8,2307.2,-11915.,25488.
566.0000000000,5435.9,2307.2,-11911.,25488.
567.0000000000,5435.9,2307.3,-11907.,25488.
568.0000000000,5436.0,2307.3,-11903.,25488.
569.0000000000,5436.0,2307.3,-11898.,25488.
570.0000000000,5436.1,2307.3,-11894.,25489.
571.0000000000,5436.1,2307.3,-11890.,25489.
572.0000000000,5436.2,2307.3,-11886.,25489.
573.0000000000,5436.3,2307.3,-11882.,25489.
574.0000000000,5436.3,2307.4,-11877.,25489.
575.0000000000,5436.4,2307.4,-11873.,25489.
576.0000000000,5436.4,2307.4,-11869.,25489.
577.0000000000,5436.5,2307.4,-11865.,25489.
578.0000000000,5436.5,2307.4,-11860.,25489.
579.0000000000,5436.6,2307.4,-11857.,25490.
580.0000000000,5436.6,2307.5,-11854.,25490.
581.0000000000,5436.7,2307.5,-11851.,25490.
582.0000000000,5436.7,2307.5,-11847.,25490.
583.0000000000,5436.8,2307.5,-11843.,25490.
584.0000000000,5436.8,2307.5,-11839.,25490.
585.0000000000,5436.9,2307.5,-11835.,25490.
586.0000000000,5437.0,2307.6,-11831.,25490.
587.0000000000,5437.0,2307.6,-11826.,25490.
588.0000000000,5437.1,2307.6,-11822.,25491.
589.0000000000,5437.1,2307.6,-11818.,25491.
590.0000000000,5437.2,2307.6,-11815.,25491.
591.0000000000,5437.2,2307.6,-11811.,25491.
592.0000000000,5437.3,2307.6,-11806.,25491.
593.0000000000,5437.3,2307.7,-11802.,25491.
594.0000000000,5437.4,2307.7,-11798.,25491.
595.0000000000,5437.4,2307.7,-11795.,25491.
596.0000000000,5437.5,2307.7,-11791.,25492.
597.0000000000,5437.5,2307.7,-11788.,25492.
598.0000000000,5437.6,2307.7,-11784.,25492.
599.0000000000,5437.7,2307.8,-11779.,25492.
600.0000000000,5437.7,2307.8,-11775.,25492.
601.0000000000,5437.8,2307.8,-11771.,25492.
602.0000000000,5437.8,2307.8,-11767.,25492.
603.0000000000,5437.9,2307.8,-11763.,25492.
604.0000000000,5437.9,2307.8,-11759.,25492.
605.0000000000,5438.0,2307.9,-11755.,25493.
606.0000000000,5438.0,2307.9,-11751.,25493.
607.0000000000,5438.1,2307.9,-11747.,25493.
608.0000000000,5438.1,2307.9,-11743.,25493.
609.0000000000,5438.2,2307.9,-11739.,25493.
610.0000000000,5438.3,2307.9,-11734.,25493.
611.0000000000,5438.3,2308.0,-11730.,25493.
612.0000000000,5438.4,2308.0,-11726.,25493.
613.0000000000,5438.4,2308.0,-11723.,25494.
614.0000000000,5438.5,2308.0,-11719.,25494.
615.0000000000,5438.5,2308.0,-11715.,25494.
616.0000000000,5438.6,2308.0,-11711.,25494.
617.0000000000,5438.6,2308.1,-11707.,25494.
618.0000000000,5438.7,2308.1,-11703.,25494.
619.0000000000,5438.7,2308.1,-11699.,25494.
620.0000000000,5438.8,2308.1,-11695.,25494.
621.0000000000,5438.9,2308.1,-11691.,25495.
622.0000000000,5438.9,2308.1,-11688.,25495.
623.0000000000,5439.0,2308.1,-11684.,25495.
624.0000000000,5439.0,2308.2,-11680.,25495.
625.0000000000,5439.1,2308.2,-11676.,25495.
626.0000000000,5439.1,2308.2,-11672.,25495.
627.0000000000,5439.2,2308.2,-11668.,25495.
628.0000000000,5439.2,2308.2,-11665.,25495.
629.0000000000,5439.3,2308.2,-11661.,25495.
630.0000000000,5439.3,2308.3,-11658.,25496.
631.0000000000,5439.4,2308.3,-11654.,25496.
632.0000000000,5439.5,2308.3,-11650.,25496.
633.0000000000,5439.5,2308.3,-11646.,25496.
634.0000000000,5439.6,2308.3,-11642.,25496.
635.0000000000,5439.6,2308.3,-11640.,25496.
636.0000000000,5439.7,2308.4,-11637.,25496.
637.0000000000,5439.7,2308.4,-11633.,25496.
638.0000000000,5439.8,2308.4,-11630.,25497.
639.0000000000,5439.8,2308.4,-11626.,25497.
640.0000000000,5439.9,2308.4,-11622.,25497.
641.0000000000,5440.0,2308.4,-11618.,25497.
642.0000000000,5440.0,2308.5,-11614.,25497.
643.0000000000,5440.1,2308.5,-11610.,25497.
644.0000000000,5440.1,2308.5,-11606.,25497.
645.0000000000,5440.2,2308.5,-11602.,25497.
646.0000000000,5440.2,2308.5,-11598.,25498.
647.0000000000,5440.3,2308.5,-11594.,25498.
648.0000000000,5440.3,2308.6,-11590.,25498.
649.0000000000,5440.4,2308.6,-11587.,25498.
650.0000000000,5440.5,2308.6,-11583.,25498.
651.0000000000,5440.5,2308.6,-11579.,25498.
652.0000000000,5440.6,2308.6,-11575.,25498.
653.0000000000,5440.6,2308.6,-11571.,25498.
654.0000000000,5440.7,2308.7,-11567.,25499.
655.0000000000,5440.7,2308.7,-11563.,25499.
656.0000000000,5440.8,2308.7,-11559.,25499.
657.0000000000,5440.8,2308.7,-11555.,25499.
658.0000000000,5440.9,2308.7,-11551.,25499.
659.0000000000,5440.9,2308.7,-11547.,25499.
660.0000000000,5441.0,2308.8,-11544.,25499.
661.0000000000,5441.1,2308.8,-11540.,25499.
662.0000000000,5441.1,2308.8,-11536.,25500.
663.0000000000,5441.2,2308.8,-11533.,25500.
664.0000000000,5441.2,2308.8,-11529.,25500.
665.0000000000,5441.3,2308.8,-11525.,25500.
666.0000000000,5441.3,2308.9,-11521.,25500.
667.0000000000,5441.4,2308.9,-11517.,25500.
668.0000000000,5441.5,2308.9,-11513.,25500.
669.0000000000,5441.5,2308.9,-11509.,25500.
670.0000000000,5441.6,2308.9,-11505.,25501.
671.0000000000,5441.6,2308.9,-11501.,25501.
672.0000000000,5441.7,2309.0,-11497.,25501.
673.0000000000,5441.7,2309.0,-11493.,25501.
674.0000000000,5441.8,2309.0,-11492.,25501.
675.0000000000,5441.8,2309.0,-11490.,25501.
676.0000000000,5441.9,2309.0,-11488.,25501.
677.0000000000,5442.0,2309.0,-11484.,25501.
678.0000000000,5442.0,2309.1,-11480.,25502.
679.0000000000,5442.1,2309.1,-11477.,25502.
680.0000000000,5442.1,2309.1,-11473.,25502.
681.0000000000,5442.2,2309.1,-11469.,25502.
682.0000000000,5442.2,2309.1,-11465.,25502.
683.0000000000,5442.3,2309.1,-11461.,25502.
684.0000000000,5442.3,2309.2,-11457.,25502.
685.0000000000,5442.4,2309.2,-11453.,25502.
686.0000000000,5442.5,2309.2,-11449.,25503.
687.0000000000,5442.5,2309.2,-11446.,25503.
688.0000000000,5442.6,2309.2,-11442.,25503.
689.0000000000,5442.6,2309.2,-11438.,25503.
690.0000000000,5442.7,2309.3,-11434.,25503.
691.0000000000,5442.7,2309.3,-11430.,25503.
692.0000000000,5442.8,2309.3,-11426.,25503.
693.0000000000,5442.9,2309.3,-11423.,25503.
694.0000000000,5442.9,2309.3,-11419.,25504.
695.0000000000,5443.0,2309.3,-11415.,25504.
696.0000000000,5443.0,2309.4,-11411.,25504.
697.0000000000,5443.1,2309.4,-11407.,25504.
698.0000000000,5443.1,2309.4,-11403.,25504.
699.0000000000,5443.2,2309.4,-11399.,25504.
700.0000000000,5443.2,2309.4,-11395.,25504.
701.0000000000,5443.3,2309.4,-11392.,25505.
702.0000000000,5443.4,2309.5,-11388.,25505.
703.0000000000,5443.4,2309.5,-11384.,25505.
704.0000000000,5443.5,2309.5,-11380.,25505.
705.0000000000,5443.5,2309.5,-11376.,25505.
706.0000000000,5443.6,2309.5,-11372.,25505.
707.0000000000,5443.6,2309.5,-11368.,25505.
708.0000000000,5443.7,2309.6,-11365.,25505.
709.0000000000,5443.8,2309.6,-11361.,25506.
710.0000000000,5443.8,2309.6,-11357.,25506.
711.0000000000,5443.9,2309.6,-11353.,25506.
712.0000000000,5443.9,2309.6,-11349.,25506.
713.0000000000,5444.0,2309.6,-11345.,25506.
714.0000000000,5444.0,2309.7,-11342.,25506.
715.0000000000,5444.1,2309.7,-11338.,25506.
716.0000000000,5444.1,2309.7,-11334.,25506.
717.0000000000,5444.2,2309.7,-11330.,25507.
718.0000000000,5444.3,2309.7,-11326.,25507.
719.0000000000,5444.3,2309.8,-11322.,25507.
720.0000000000,5444.4,2309.8,-11319.,25507.
721.0000000000,5444.4,2309.8,-11315.,25507.
722.0000000000,5444.5,2309.8,-11311.,25507.
723.0000000000,5444.5,2309.8,-11307.,25507.
724.0000000000,5444.6,2309.8,-11303.,25508.
725.0000000000,5444.7,2309.9,-11299.,25508.
726.0000000000,5444.7,2309.9,-11296.,25508.
727.0000000000,5444.8,2309.9,-11293.,25508.
728.0000000000,5444.8,2309.9,-11289.,25508.
729.0000000000,5444.9,2309.9,-11286.,25508.
730.0000000000,5444.9,2309.9,-11282.,25508.
731.0000000000,5445.0,2310.0,-11279.,25508.
732.0000000000,5445.1,2310.0,-11275.,25509.
733.0000000000,5445.1,2310.0,-11272.,25509.
734.0000000000,5445.2,2310.0,-11268.,25509.
735.0000000000,5445.2,2310.0,-11265.,25509.
736.0000000000,5445.3,2310.0,-11261.,25509.
737.0000000000,5445.3,2310.1,-11257.,25509.
738.0000000000,5445.4,2310.1,-11253.,25509.
739.0000000000,5445.4,2310.1,-11249.,25509.
740.0000000000,5445.4,2310.1,-11246.,25510.
741.0000000000,5445.5,2310.1,-11242.,25510.
742.0000000000,5445.5,2310.1,-11239.,25510.
743.0000000000,5445.6,2310.2,-11235.,25510.
744.0000000000,5445.6,2310.2,-11231.,25510.
745.0000000000,5445.7,2310.2,-11227.,25510.
746.0000000000,5445.7,2310.2,-11224.,25510.
747.0000000000,5445.8,2310.2,-11220.,25511.
748.0000000000,5445.8,2310.3,-11216.,25511.
749.0000000000,5445.9,2310.3,-11212.,25511.
750.0000000000,5445.9,2310.3,-11208.,25511.
751.0000000000,5446.0,2310.3,-11205.,25511.
752.0000000000,5446.0,2310.3,-11201.,25511.
753.0000000000,5446.1,2310.3,-11198.,25511.
754.0000000000,5446.2,2310.3,-11194.,25511.
755.0000000000,5446.2,2310.3,-11191.,25512.
756.0000000000,5446.3,2310.3,-11187.,25512.
757.0000000000,5446.3,2310.3,-11183.,25512.
758.0000000000,5446.4,2310.3,-11179.,25512.
759.0000000000,5446.4,2310.3,-11176.,25512.
760.0000000000,5446.5,2310.3,-11172.,25512.
761.0000000000,5446.6,2310.3,-11168.,25512.
762.0000000000,5446.6,2310.3,-11165.,25513.
763.0000000000,5446.7,2310.3,-11162.,25513.
764.0000000000,5446.7,2310.3,-11158.,25513.
765.0000000000,5446.8,2310.3,-11154.,25513.
766.0000000000,5446.8,2310.3,-11150.,25513.
767.0000000000,5446.9,2310.3,-11147.,25513.
768.0000000000,5447.0,2310.3,-11143.,25513.
769.0000000000,5447.0,2310.3,-11139.,25513.
770.0000000000,5447.1,2310.4,-11135.,25514.
771.0000000000,5447.1,2310.4,-11132.,25514.
772.0000000000,5447.2,2310.4,-11128.,25514.
773.0000000000,5447.2,2310.4,-11124.,25514.
774.0000000000,5447.3,2310.4,-11120.,25514.
775.0000000000,5447.4,2310.4,-11117.,25514.
776.0000000000,5447.4,2310.4,-11113.,25514.
777.0000000000,5447.5,2310.4,-11109.,25515.
778.0000000000,5447.5,2310.5,-11105.,25515.
779.0000000000,5447.6,2310.5,-11102.,25515.
780.0000000000,5447.6,2310.5,-11098.,25515.
781.0000000000,5447.7,2310.5,-11094.,25515.
782.0000000000,5447.8,2310.5,-11091.,25515.
783.0000000000,5447.8,2310.5,-11087.,25515.
784.0000000000,5447.9,2310.6,-11083.,25516.
785.0000000000,5447.9,2310.6,-11079.,25516.
786.0000000000,5448.0,2310.6,-11076.,25516.
787.0000000000,5448.0,2310.6,-11072.,25516.
788.0000000000,5448.1,2310.6,-11068.,25516.
789.0000000000,5448.2,2310.6,-11064.,25516.
790.0000000000,5448.2,2310.7,-11061.,25516.
791.0000000000,5448.3,2310.7,-11057.,25516.
792.0000000000,5448.3,2310.7,-11053.,25517.
793.0000000000,5448.4,2310.7,-11050.,25517.
794.0000000000,5448.4,2310.7,-11047.,25517.
795.0000000000,5448.5,2310.7,-11043.,25517.
796.0000000000,5448.6,2310.8,-11039.,25517.
797.0000000000,5448.6,2310.8,-11036.,25517.
798.0000000000,5448.7,2310.8,-11032.,25517.
799.0000000000,5448.7,2310.8,-11029.,25518.
800.0000000000,5448.8,2310.8,-11025.,25518.
801.0000000000,5448.9,2310.9,-11021.,25518.
802.0000000000,5448.9,2310.9,-11018.,25518.
803.0000000000,5449.0,2310.9,-11014.,25518.
804.0000000000,5449.0,2310.9,-11010.,25518.
805.0000000000,5449.1,2310.9,-11007.,25518.
806.0000000000,5449.1,2310.9,-11003.,25519.
807.0000000000,5449.2,2311.0,-10999.,25519.
808.0000000000,5449.3,2311.0,-10996.,25519.
809.0000000000,5449.3,2311.0,-10993.,25519.
810.0000000000,5449.4,2311.0,-10991.,25519.
811.0000000000,5449.4,2311.0,-10989.,25519.
812.0000000000,5449.5,2311.0,-10986.,25519.
813.0000000000,5449.5,2311.1,-10983.,25520.
814.0000000000,5449.6,2311.1,-10980.,25520.
815.0000000000,5449.7,2311.1,-10976.,25520.
816.0000000000,5449.7,2311.1,-10972.,25520.
817.0000000000,5449.8,2311.1,-10969.,25520.
818.0000000000,5449.8,2311.2,-10965.,25520.
819.0000000000,5449.9,2311.2,-10962.,25520.
820.0000000000,5450.0,2311.2,-10958.,25520.
821.0000000000,5450.0,2311.2,-10954.,25521.
822.0000000000,5450.1,2311.2,-10951.,25521.
823.0000000000,5450.1,2311.2,-10947.,25521.
824.0000000000,5450.2,2311.3,-10943.,25521.
825.0000000000,5450.2,2311.3,-10940.,25521.
826.0000000000,5450.3,2311.3,-10936.,25521.
827.0000000000,5450.4,2311.3,-10933.,25521.
828.0000000000,5450.4,2311.3,-10929.,25522.
829.0000000000,5450.5,2311.4,-10926.,25522.
830.0000000000,5450.5,2311.4,-10922.,25522.
831.0000000000,5450.6,2311.4,-10919.,25522.
832.0000000000,5450.7,2311.4,-10915.,25522.
833.0000000000,5450.7,2311.4,-10912.,25522.
834.0000000000,5450.8,2311.5,-10909.,25522.
835.0000000000,5450.8,2311.5,-10906.,25523.
836.0000000000,5450.9,2311.5,-10903.,25523.
837.0000000000,5450.9,2311.5,-10899.,25523.
838.0000000000,5451.0,2311.5,-10897.,25523.
839.0000000000,5451.1,2311.5,-10893.,25523.
840.0000000000,5451.1,2311.6,-10890.,25523.
841.0000000000,5451.2,2311.6,-10886.,25523.
842.0000000000,5451.2,2311.6,-10883.,25524.
843.0000000000,5451.3,2311.6,-10879.,25524.
844.0000000000,5451.4,2311.6,-10876.,25524.
845.0000000000,5451.4,2311.7,-10873.,25524.
846.0000000000,5451.5,2311.7,-10869.,25524.
847.0000000000,5451.5,2311.7,-10866.,25524.
848.0000000000,5451.6,2311.7,-10863.,25524.
849.0000000000,5451.7,2311.7,-10860.,25524.
850.0000000000,5451.7,2311.8,-10856.,25525.
851.0000000000,5451.8,2311.8,-10853.,25525.
852.0000000000,5451.8,2311.8,-10849.,25525.
853.0000000000,5451.9,2311.8,-10846.,25525.
854.0000000000,5451.9,2311.8,-10842.,25525.
855.0000000000,5452.0,2311.8,-10839.,25525.
856.0000000000,5452.1,2311.9,-10835.,25525.
857.0000000000,5452.1,2311.9,-10832.,25526.
858.0000000000,5452.2,2311.9,-10828.,25526.
859.0000000000,5452.2,2311.9,-10825.,25526.
860.0000000000,5452.3,2311.9,-10821.,25526.
861.0000000000,5452.4,2312.0,-10820.,25526.
862.0000000000,5452.4,2312.0,-10819.,25526.
863.0000000000,5452.5,2312.0,-10818.,25526.
864.0000000000,5452.5,2312.0,-10816.,25527.
865.0000000000,5452.6,2312.0,-10813.,25527.
866.0000000000,5452.7,2312.1,-10811.,25527.
867.0000000000,5452.7,2312.1,-10810.,25527.
868.0000000000,5452.8,2312.1,-10808.,25527.
869.0000000000,5452.8,2312.1,-10805.,25527.
870.0000000000,5452.9,2312.1,-10801.,25527.
871.0000000000,5452.9,2312.1,-10799.,25528.
872.0000000000,5453.0,2312.2,-10796.,25528.
873.0000000000,5453.1,2312.2,-10793.,25528.
874.0000000000,5453.1,2312.2,-10790.,25528.
875.0000000000,5453.2,2312.2,-10787.,25528.
876.0000000000,5453.2,2312.2,-10783.,25528.
877.0000000000,5453.3,2312.3,-10780.,25528.
878.0000000000,5453.4,2312.3,-10777.,25528.
879.0000000000,5453.4,2312.3,-10775.,25529.
880.0000000000,5453.5,2312.3,-10773.,25529.
881.0000000000,5453.5,2312.3,-10771.,25529.
882.0000000000,5453.6,2312.4,-10768.,25529.
883.0000000000,5453.7,2312.4,-10765.,25529.
884.0000000000,5453.7,2312.4,-10762.,25529.
885.0000000000,5453.8,2312.4,-10759.,25529.
886.0000000000,5453.8,2312.4,-10755.,25530.
887.0000000000,5453.9,2312.4,-10752.,25530.
888.0000000000,5453.9,2312.5,-10748.,25530.
889.0000000000,5454.0,2312.5,-10745.,25530.
890.0000000000,5454.1,2312.5,-10741.,25530.
891.0000000000,5454.1,2312.5,-10738.,25530.
892.0000000000,5454.2,2312.5,-10735.,25530.
893.0000000000,5454.2,2312.6,-10731.,25531.
894.0000000000,5454.3,2312.6,-10728.,25531.
895.0000000000,5454.3,2312.6,-10726.,25531.
896.0000000000,5454.4,2312.6,-10723.,25531.
897.0000000000,5454.5,2312.6,-10720.,25531.
898.0000000000,5454.5,2312.7,-10718.,25531.
899.0000000000,5454.6,2312.7,-10715.,25531.
900.0000000000,5454.6,2312.7,-10711.,25532.
901.0000000000,5454.7,2312.7,-10709.,25532.
902.0000000000,5454.8,2312.7,-10705.,25532.
903.0000000000,5454.8,2312.8,-10702.,25532.
904.0000000000,5454.9,2312.8,-10699.,25532.
905.0000000000,5454.9,2312.8,-10696.,25532.
906.0000000000,5455.0,2312.8,-10692.,25532.
907.0000000000,5455.0,2312.8,-10689.,25533.
908.0000000000,5455.1,2312.8,-10686.,25533.
909.0000000000,5455.2,2312.9,-10684.,25533.
910.0000000000,5455.2,2312.9,-10681.,25533.
911.0000000000,5455.3,2312.9,-10678.,25533.
912.0000000000,5455.3,2312.9,-10674.,25533.
913.0000000000,5455.4,2312.9,-10671.,25533.
914.0000000000,5455.5,2313.0,-10668.,25534.
915.0000000000,5455.5,2313.0,-10664.,25534.
916.0000000000,5455.6,2313.0,-10661.,25534.
917.0000000000,5455.6,2313.0,-10658.,25534.
918.0000000000,5455.7,2313.0,-10654.,25534.
919.0000000000,5455.7,2313.1,-10652.,25534.
920.0000000000,5455.8,2313.1,-10648.,25534.
921.0000000000,5455.9,2313.1,-10645.,25534.
922.0000000000,5455.9,2313.1,-10642.,25535.
923.0000000000,5456.0,2313.1,-10638.,25535.
924.0000000000,5456.0,2313.2,-10635.,25535.
925.0000000000,5456.1,2313.2,-10632.,25535.
926.0000000000,5456.2,2313.2,-10628.,25535.
927.0000000000,5456.2,2313.2,-10625.,25535.
928.0000000000,5456.3,2313.2,-10621.,25535.
929.0000000000,5456.3,2313.2,-10618.,25536.
930.0000000000,5456.4,2313.3,-10615.,25536.
931.0000000000,5456.4,2313.3,-10611.,25536.
932.0000000000,5456.5,2313.3,-10608.,25536.
933.0000000000,5456.6,2313.3,-10604.,25536.
934.0000000000,5456.6,2313.3,-10601.,25536.
935.0000000000,5456.7,2313.4,-10598.,25536.
936.0000000000,5456.7,2313.4,-10594.,25537.
937.0000000000,5456.8,2313.4,-10591.,25537.
938.0000000000,5456.9,2313.4,-10587.,25537.
939.0000000000,5456.9,2313.4,-10584.,25537.
940.0000000000,5457.0,2313.5,-10581.,25537.
941.0000000000,5457.0,2313.5,-10577.,25537.
942.0000000000,5457.1,2313.5,-10574.,25537.
943.0000000000,5457.1,2313.5,-10571.,25538.
944.0000000000,5457.2,2313.5,-10568.,25538.
945.0000000000,5457.3,2313.6,-10564.,25538.
946.0000000000,5457.3,2313.6,-10561.,25538.
947.0000000000,5457.4,2313.6,-10558.,25538.
948.0000000000,5457.4,2313.6,-10554.,25538.
949.0000000000,5457.5,2313.6,-10551.,25538.
950.0000000000,5457.6,2313.7,-10548.,25539.
951.0000000000,5457.6,2313.7,-10544.,25539.
952.0000000000,5457.7,2313.7,-10541.,25539.
953.0000000000,5457.7,2313.7,-10537.,25539.
954.0000000000,5457.8,2313.7,-10534.,25539.
955.0000000000,5457.8,2313.8,-10531.,25539.
956.0000000000,5457.9,2313.8,-10528.,25539.
957.0000000000,5458.0,2313.8,-10525.,25540.
958.0000000000,5458.0,2313.8,-10522.,25540.
959.0000000000,5458.1,2313.8,-10519.,25540.
960.0000000000,5458.1,2313.8,-10516.,25540.
961.0000000000,5458.2,2313.9,-10513.,25540.
962.0000000000,5458.3,2313.9,-10510.,25540.
963.0000000000,5458.3,2313.9,-10507.,25540.
964.0000000000,5458.4,2313.9,-10504.,25541.
965.0000000000,5458.4,2313.9,-10501.,25541.
966.0000000000,5458.5,2314.0,-10498.,25541.
967.0000000000,5458.6,2314.0,-10494.,25541.
968.0000000000,5458.6,2314.0,-10491.,25541.
969.0000000000,5458.7,2314.0,-10488.,25541.
970.0000000000,5458.7,2314.0,-10485.,25541.
971.0000000000,5458.8,2314.1,-10482.,25542.
972.0000000000,5458.9,2314.1,-10478.,25542.
973.0000000000,5458.9,2314.1,-10475.,25542.
974.0000000000,5459.0,2314.1,-10472.,25542.
975.0000000000,5459.0,2314.1,-10468.,25542.
976.0000000000,5459.1,2314.2,-10465.,25542.
977.0000000000,5459.1,2314.2,-10462.,25542.
978.0000000000,5459.2,2314.2,-10459.,25543.
979.0000000000,5459.3,2314.2,-10455.,25543.
980.0000000000,5459.3,2314.2,-10452.,25543.
981.0000000000,5459.4,2314.3,-10449.,25543.
982.0000000000,5459.4,2314.3,-10445.,25543.
983.0000000000,5459.5,2314.3,-10442.,25543.
984.0000000000,5459.6,2314.3,-10439.,25543.
985.0000000000,5459.6,2314.3,-10436.,25544.
986.0000000000,5459.7,2314.4,-10433.,25544.
987.0000000000,5459.7,2314.4,-10430.,25544.
988.0000000000,5459.8,2314.4,-10426.,25544.
989.0000000000,5459.9,2314.4,-10423.,25544.
990.0000000000,5459.9,2314.4,-10420.,25544.
991.0000000000,5460.0,2314.5,-10417.,25544.
992.0000000000,5460.0,2314.5,-10413.,25545.
993.0000000000,5460.1,2314.5,-10410.,25545.
994.0000000000,5460.2,2314.5,-10407.,25545.
995.0000000000,5460.2,2314.5,-10403.,25545.
996.0000000000,5460.3,2314.6,-10400.,25545.
997.0000000000,5460.3,2314.6,-10397.,25545.
998.0000000000,5460.4,2314.6,-10393.,25545.
999.0000000000,5460.5,2314.6,-10390.,25546.
1000.000000000,5460.5,2314.6,-10387.,25546.
1001.000000000,5460.6,2314.7,-10384.,25546.
1002.000000000,5460.6,2314.7,-10381.,25546.
1003.000000000,5460.7,2314.7,-10377.,25546.
1004.000000000,5460.8,2314.7,-10374.,25546.
1005.000000000,5460.8,2314.7,-10371.,25546.
1006.000000000,5460.9,2314.8,-10367.,25547.
1007.000000000,5460.9,2314.8,-10364.,25547.
1008.000000000,5461.0,2314.8,-10361.,25547.
1009.000000000,5461.1,2314.8,-10358.,25547.
1010.000000000,5461.1,2314.8,-10354.,25547.
1011.000000000,5461.2,2314.9,-10351.,25547.
1012.000000000,5461.2,2314.9,-10350.,25547.
1013.000000000,5461.3,2314.9,-10347.,25548.
1014.000000000,5461.4,2314.9,-10345.,25548.
1015.000000000,5461.4,2314.9,-10342.,25548.
1016.000000000,5461.5,2315.0,-10339.,25548.
1017.000000000,5461.5,2315.0,-10335.,25548.
1018.000000000,5461.6,2315.0,-10332.,25548.
1019.000000000,5461.7,2315.0,-10329.,25548.
1020.000000000,5461.7,2315.0,-10326.,25549.
1021.000000000,5461.8,2315.1,-10322.,25549.
1022.000000000,5461.8,2315.1,-10319.,25549.
1023.000000000,5461.9,2315.1,-10316.,25549.
1024.000000000,5462.0,2315.1,-10313.,25549.
1025.000000000,5462.0,2315.1,-10309.,25549.
1026.000000000,5462.1,2315.2,-10306.,25549.
1027.000000000,5462.1,2315.2,-10307.,25550.
1028.000000000,5462.2,2315.2,-10307.,25550.
1029.000000000,5462.3,2315.2,-10305.,25550.
1030.000000000,5462.3,2315.2,-10303.,25550.
1031.000000000,5462.4,2315.3,-10300.,25550.
1032.000000000,5462.4,2315.3,-10297.,25550.
1033.000000000,5462.5,2315.3,-10294.,25550.
1034.000000000,5462.6,2315.3,-10293.,25551.
1035.000000000,5462.6,2315.3,-10291.,25551.
1036.000000000,5462.7,2315.4,-10288.,25551.
1037.000000000,5462.7,2315.4,-10285.,25551.
1038.000000000,5462.8,2315.4,-10282.,25551.
1039.000000000,5462.9,2315.4,-10279.,25551.
1040.000000000,5462.9,2315.4,-10276.,25551.
1041.000000000,5463.0,2315.5,-10272.,25552.
1042.000000000,5463.0,2315.5,-10269.,25552.
1043.000000000,5463.1,2315.5,-10266.,25552.
1044.000000000,5463.2,2315.5,-10263.,25552.
1045.000000000,5463.2,2315.5,-10260.,25552.
1046.000000000,5463.3,2315.6,-10257.,25552.
1047.000000000,5463.3,2315.6,-10253.,25552.
1048.000000000,5463.4,2315.6,-10250.,25553.
1049.000000000,5463.5,2315.6,-10247.,25553.
1050.000000000,5463.5,2315.6,-10244.,25553.
1051.000000000,5463.6,2315.7,-10241.,25553.
1052.000000000,5463.7,2315.7,-10238.,25553.
1053.000000000,5463.7,2315.7,-10235.,25553.
1054.000000000,5463.8,2315.7,-10231.,25553.
1055.000000000,5463.8,2315.7,-10228.,25554.
1056.000000000,5463.9,2315.8,-10225.,25554.
1057.000000000,5464.0,2315.8,-10222.,25554.
1058.000000000,5464.0,2315.8,-10219.,25554.
1059.000000000,5464.1,2315.8,-10215.,25554.
1060.000000000,5464.1,2315.8,-10212.,25554.
1061.000000000,5464.2,2315.9,-10209.,25554.
1062.000000000,5464.3,2315.9,-10208.,25555.
1063.000000000,5464.3,2315.9,-10205.,25555.
1064.000000000,5464.4,2315.9,-10202.,25555.
1065.000000000,5464.4,2315.9,-10199.,25555.
1066.000000000,5464.5,2316.0,-10196.,25555.
1067.000000000,5464.6,2316.0,-10193.,25555.
1068.000000000,5464.6,2316.0,-10190.,25555.
1069.000000000,5464.7,2316.0,-10187.,25556.
1070.000000000,5464.7,2316.0,-10183.,25556.
1071.000000000,5464.8,2316.1,-10180.,25556.
1072.000000000,5464.9,2316.1,-10177.,25556.
1073.000000000,5464.9,2316.1,-10174.,25556.
1074.000000000,5465.0,2316.1,-10171.,25556.
1075.000000000,5465.0,2316.1,-10167.,25557.
1076.000000000,5465.1,2316.2,-10164.,25557.
1077.000000000,5465.2,2316.2,-10163.,25557.
1078.000000000,5465.2,2316.2,-10160.,25557.
1079.000000000,5465.3,2316.2,-10157.,25557.
1080.000000000,5465.3,2316.2,-10154.,25557.
1081.000000000,5465.4,2316.3,-10151.,25557.
1082.000000000,5465.5,2316.3,-10148.,25558.
1083.000000000,5465.5,2316.3,-10145.,25558.
1084.000000000,5465.6,2316.3,-10142.,25558.
1085.000000000,5465.6,2316.3,-10138.,25558.
1086.000000000,5465.7,2316.4,-10135.,25558.
1087.000000000,5465.8,2316.4,-10132.,25558.
1088.000000000,5465.8,2316.4,-10129.,25558.
1089.000000000,5465.9,2316.4,-10126.,25559.
1090.000000000,5465.9,2316.4,-10123.,25559.
1091.000000000,5466.0,2316.5,-10121.,25559.
1092.000000000,5466.1,2316.5,-10118.,25559.
1093.000000000,5466.1,2316.5,-10116.,25559.
1094.000000000,5466.2,2316.5,-10113.,25559.
1095.000000000,5466.2,2316.5,-10110.,25559.
1096.000000000,5466.3,2316.6,-10106.,25560.
1097.000000000,5466.4,2316.6,-10103.,25560.
1098.000000000,5466.4,2316.6,-10100.,25560.
1099.000000000,5466.5,2316.6,-10097.,25560.
1100.000000000,5466.5,2316.6,-10094.,25560.
1101.000000000,5466.6,2316.7,-10091.,25560.
1102.000000000,5466.7,2316.7,-10088.,25560.
1103.000000000,5466.7,2316.7,-10085.,25561.
1104.000000000,5466.8,2316.7,-10082.,25561.
1105.000000000,5466.9,2316.8,-10079.,25561.
1106.000000000,5466.9,2316.8,-10075.,25561.
1107.000000000,5467.0,2316.8,-10072.,25561.
1108.000000000,5467.0,2316.8,-10069.,25561.
1109.000000000,5467.1,2316.8,-10066.,25561.
1110.000000000,5467.2,2316.9,-10063.,25562.
1111.000000000,5467.2,2316.9,-10060.,25562.
1112.000000000,5467.3,2316.9,-10057.,25562.
1113.000000000,5467.3,2316.9,-10053.,25562.
1114.000000000,5467.4,2316.9,-10050.,25562.
1115.000000000,5467.5,2317.0,-10047.,25562.
1116.000000000,5467.5,2317.0,-10044.,25562.
1117.000000000,5467.6,2317.0,-10041.,25563.
1118.000000000,5467.6,2317.0,-10038.,25563.
1119.000000000,5467.7,2317.0,-10035.,25563.
1120.000000000,5467.8,2317.1,-10032.,25563.
1121.000000000,5467.8,2317.1,-10028.,25563.
1122.000000000,5467.9,2317.1,-10026.,25563.
1123.000000000,5468.0,2317.1,-10023.,25563.
1124.000000000,5468.0,2317.1,-10020.,25564.
1125.000000000,5468.1,2317.2,-10017.,25564.
1126.000000000,5468.1,2317.2,-10014.,25564.
1127.000000000,5468.2,2317.2,-10011.,25564.
1128.000000000,5468.3,2317.2,-10008.,25564.
1129.000000000,5468.3,2317.2,-10005.,25564.
1130.000000000,5468.4,2317.3,-10002.,25564.
1131.000000000,5468.4,2317.3,-9998.8,25565.
1132.000000000,5468.5,2317.3,-9995.7,25565.
1133.000000000,5468.6,2317.3,-9992.6,25565.
1134.000000000,5468.6,2317.3,-9989.5,25565.
1135.000000000,5468.7,2317.4,-9986.4,25565.
1136.000000000,5468.7,2317.4,-9983.3,25565.
1137.000000000,5468.8,2317.4,-9980.2,25566.
1138.000000000,5468.9,2317.4,-9977.1,25566.
1139.000000000,5468.9,2317.5,-9974.0,25566.
1140.000000000,5469.0,2317.5,-9970.9,25566.
1141.000000000,5469.1,2317.5,-9967.8,25566.
1142.000000000,5469.1,2317.5,-9964.7,25566.
1143.000000000,5469.2,2317.5,-9961.7,25566.
1144.000000000,5469.2,2317.6,-9958.6,25567.
1145.000000000,5469.3,2317.6,-9955.5,25567.
1146.000000000,5469.4,2317.6,-9952.4,25567.
1147.000000000,5469.4,2317.6,-9949.4,25567.
1148.000000000,5469.5,2317.6,-9946.6,25567.
1149.000000000,5469.6,2317.7,-9944.6,25567.
1150.000000000,5469.6,2317.7,-9941.9,25567.
1151.000000000,5469.7,2317.7,-9939.1,25568.
1152.000000000,5469.7,2317.7,-9936.1,25568.
1153.000000000,5469.8,2317.7,-9933.1,25568.
1154.000000000,5469.9,2317.8,-9930.0,25568.
1155.000000000,5469.9,2317.8,-9927.0,25568.
1156.000000000,5470.0,2317.8,-9923.9,25568.
1157.000000000,5470.0,2317.8,-9920.9,25568.
1158.000000000,5470.1,2317.8,-9917.8,25569.
1159.000000000,5470.2,2317.9,-9914.7,25569.
1160.000000000,5470.2,2317.9,-9911.7,25569.
1161.000000000,5470.3,2317.9,-9908.6,25569.
1162.000000000,5470.4,2317.9,-9905.6,25569.
1163.000000000,5470.4,2318.0,-9904.0,25569.
1164.000000000,5470.5,2318.0,-9902.6,25569.
1165.000000000,5470.5,2318.0,-9901.6,25570.
1166.000000000,5470.6,2318.0,-9900.9,25570.
1167.000000000,5470.7,2318.0,-9899.7,25570.
1168.000000000,5470.7,2318.1,-9897.5,25570.
1169.000000000,5470.8,2318.1,-9894.9,25570.
1170.000000000,5470.9,2318.1,-9892.0,25570.
1171.000000000,5470.9,2318.1,-9889.1,25571.
1172.000000000,5471.0,2318.1,-9886.1,25571.
1173.000000000,5471.0,2318.2,-9883.1,25571.
1174.000000000,5471.1,2318.2,-9880.8,25571.
1175.000000000,5471.2,2318.2,-9878.1,25571.
1176.000000000,5471.2,2318.2,-9875.2,25571.
1177.000000000,5471.3,2318.2,-9872.3,25571.
1178.000000000,5471.4,2318.3,-9869.3,25572.
1179.000000000,5471.4,2318.3,-9866.3,25572.
1180.000000000,5471.5,2318.3,-9863.4,25572.
1181.000000000,5471.5,2318.3,-9860.4,25572.
1182.000000000,5471.6,2318.3,-9857.4,25572.
1183.000000000,5471.7,2318.4,-9854.4,25572.
1184.000000000,5471.7,2318.4,-9851.4,25572.
1185.000000000,5471.8,2318.4,-9848.3,25573.
1186.000000000,5471.9,2318.4,-9845.3,25573.
1187.000000000,5471.9,2318.5,-9842.3,25573.
1188.000000000,5472.0,2318.5,-9839.3,25573.
1189.000000000,5472.0,2318.5,-9836.3,25573.
1190.000000000,5472.1,2318.5,-9833.3,25573.
1191.000000000,5472.2,2318.5,-9830.3,25573.
1192.000000000,5472.2,2318.6,-9827.3,25574.
1193.000000000,5472.3,2318.6,-9824.3,25574.
1194.000000000,5472.3,2318.6,-9821.3,25574.
1195.000000000,5472.4,2318.6,-9818.2,25574.
1196.000000000,5472.5,2318.6,-9815.1,25574.
1197.000000000,5472.5,2318.7,-9812.0,25574.
1198.000000000,5472.6,2318.7,-9808.9,25574.
1199.000000000,5472.7,2318.7,-9806.4,25575.
1200.000000000,5472.7,2318.7,-9803.6,25575.
1201.000000000,5472.8,2318.7,-9800.7,25575.
1202.000000000,5472.8,2318.8,-9797.6,25575.
1203.000000000,5472.9,2318.8,-9798.6,25575.
1204.000000000,5473.0,2318.8,-9798.3,25575.
1205.000000000,5473.0,2318.8,-9796.4,25576.
1206.000000000,5473.1,2318.9,-9793.9,25576.
1207.000000000,5473.2,2318.9,-9791.2,25576.
1208.000000000,5473.2,2318.9,-9788.3,25576.
1209.000000000,5473.3,2318.9,-9785.3,25576.
1210.000000000,5473.3,2318.9,-9782.4,25576.
1211.000000000,5473.4,2319.0,-9779.4,25576.
1212.000000000,5473.5,2319.0,-9776.4,25577.
1213.000000000,5473.5,2319.0,-9773.8,25577.
1214.000000000,5473.6,2319.0,-9771.0,25577.
1215.000000000,5473.7,2319.0,-9768.1,25577.
1216.000000000,5473.7,2319.1,-9765.1,25577.
1217.000000000,5473.8,2319.1,-9762.1,25577.
1218.000000000,5473.8,2319.1,-9759.1,25577.
1219.000000000,5473.9,2319.1,-9756.2,25578.
1220.000000000,5474.0,2319.2,-9753.2,25578.
1221.000000000,5474.0,2319.2,-9750.2,25578.
1222.000000000,5474.1,2319.2,-9747.2,25578.
1223.000000000,5474.2,2319.2,-9744.2,25578.
1224.000000000,5474.2,2319.2,-9741.3,25578.
1225.000000000,5474.3,2319.3,-9738.4,25578.
1226.000000000,5474.3,2319.3,-9735.5,25579.
1227.000000000,5474.4,2319.3,-9732.6,25579.
1228.000000000,5474.5,2319.3,-9729.6,25579.
1229.000000000,5474.5,2319.3,-9726.6,25579.
1230.000000000,5474.6,2319.4,-9723.7,25579.
1231.000000000,5474.7,2319.4,-9720.9,25579.
1232.000000000,5474.7,2319.4,-9718.2,25579.
1233.000000000,5474.8,2319.4,-9715.4,25580.
1234.000000000,5474.8,2319.5,-9712.9,25580.
1235.000000000,5474.9,2319.5,-9711.5,25580.
1236.000000000,5475.0,2319.5,-9709.5,25580.
1237.000000000,5475.0,2319.5,-9706.9,25580.
1238.000000000,5475.1,2319.5,-9704.2,25580.
1239.000000000,5475.2,2319.6,-9701.3,25581.
1240.000000000,5475.2,2319.6,-9698.4,25581.
1241.000000000,5475.3,2319.6,-9695.5,25581.
1242.000000000,5475.3,2319.6,-9692.6,25581.
1243.000000000,5475.4,2319.6,-9689.7,25581.
1244.000000000,5475.5,2319.7,-9686.7,25581.
1245.000000000,5475.5,2319.7,-9683.8,25581.
1246.000000000,5475.6,2319.7,-9680.9,25582.
1247.000000000,5475.7,2319.7,-9678.0,25582.
1248.000000000,5475.7,2319.7,-9675.3,25582.
1249.000000000,5475.8,2319.8,-9675.1,25582.
1250.000000000,5475.8,2319.8,-9673.9,25582.
1251.000000000,5475.9,2319.8,-9671.8,25582.
1252.000000000,5476.0,2319.8,-9669.3,25582.
1253.000000000,5476.0,2319.9,-9666.5,25583.
1254.000000000,5476.1,2319.9,-9663.7,25583.
1255.000000000,5476.2,2319.9,-9660.8,25583.
1256.000000000,5476.2,2319.9,-9658.0,25583.
1257.000000000,5476.3,2319.9,-9655.1,25583.
1258.000000000,5476.3,2320.0,-9652.2,25583.
1259.000000000,5476.4,2320.0,-9649.3,25583.
1260.000000000,5476.5,2320.0,-9646.4,25584.
1261.000000000,5476.5,2320.0,-9643.5,25584.
1262.000000000,5476.6,2320.0,-9640.6,25584.
1263.000000000,5476.7,2320.1,-9637.7,25584.
1264.000000000,5476.7,2320.1,-9634.8,25584.
1265.000000000,5476.8,2320.1,-9631.9,25584.
1266.000000000,5476.8,2320.1,-9629.1,25584.
1267.000000000,5476.9,2320.2,-9626.8,25585.
1268.000000000,5477.0,2320.2,-9624.1,25585.
1269.000000000,5477.0,2320.2,-9621.4,25585.
1270.000000000,5477.1,2320.2,-9618.5,25585.
1271.000000000,5477.2,2320.2,-9615.7,25585.
1272.000000000,5477.2,2320.3,-9612.8,25585.
1273.000000000,5477.3,2320.3,-9610.5,25585.
1274.000000000,5477.3,2320.3,-9612.3,25586.
1275.000000000,5477.4,2320.3,-9611.7,25586.
1276.000000000,5477.5,2320.4,-9609.8,25586.
1277.000000000,5477.5,2320.4,-9607.4,25586.
1278.000000000,5477.6,2320.4,-9604.8,25586.
1279.000000000,5477.7,2320.4,-9602.1,25586.
1280.000000000,5477.7,2320.4,-9599.3,25586.
1281.000000000,5477.8,2320.5,-9596.4,25587.
1282.000000000,5477.9,2320.5,-9593.6,25587.
1283.000000000,5477.9,2320.5,-9590.8,25587.
1284.000000000,5478.0,2320.5,-9587.9,25587.
1285.000000000,5478.0,2320.5,-9585.1,25587.
1286.000000000,5478.1,2320.6,-9582.2,25587.
1287.000000000,5478.2,2320.6,-9579.4,25587.
1288.000000000,5478.2,2320.6,-9576.6,25588.
1289.000000000,5478.3,2320.6,-9573.7,25588.
1290.000000000,5478.4,2320.7,-9570.9,25588.
1291.000000000,5478.4,2320.7,-9568.0,25588.
1292.000000000,5478.5,2320.7,-9565.2,25588.
1293.000000000,5478.5,2320.7,-9562.3,25588.
1294.000000000,5478.6,2320.7,-9559.5,25589.
1295.000000000,5478.7,2320.8,-9556.7,25589.
1296.000000000,5478.7,2320.8,-9553.8,25589.
1297.000000000,5478.8,2320.8,-9551.0,25589.
1298.000000000,5478.9,2320.8,-9548.1,25589.
1299.000000000,5478.9,2320.8,-9545.3,25589.
1300.000000000,5479.0,2320.9,-9542.5,25589.
1301.000000000,5479.1,2320.9,-9539.6,25590.
1302.000000000,5479.1,2320.9,-9536.8,25590.
1303.000000000,5479.2,2320.9,-9534.0,25590.
1304.000000000,5479.2,2321.0,-9531.6,25590.
1305.000000000,5479.3,2321.0,-9529.1,25590.
1306.000000000,5479.4,2321.0,-9526.3,25590.
1307.000000000,5479.4,2321.0,-9523.6,25590.
1308.000000000,5479.5,2321.0,-9520.8,25591.
1309.000000000,5479.6,2321.1,-9518.0,25591.
1310.000000000,5479.6,2321.1,-9515.2,25591.
1311.000000000,5479.7,2321.1,-9512.3,25591.
1312.000000000,5479.8,2321.1,-9509.5,25591.
1313.000000000,5479.8,2321.2,-9506.7,25591.
1314.000000000,5479.9,2321.2,-9503.9,25591.
1315.000000000,5479.9,2321.2,-9501.1,25592.
1316.000000000,5480.0,2321.2,-9498.2,25592.
1317.000000000,5480.1,2321.2,-9495.4,25592.
1318.000000000,5480.1,2321.3,-9492.6,25592.
1319.000000000,5480.2,2321.3,-9489.8,25592.
1320.000000000,5480.3,2321.3,-9487.0,25592.
1321.000000000,5480.3,2321.3,-9485.8,25593.
1322.000000000,5480.4,2321.4,-9485.1,25593.
1323.000000000,5480.5,2321.4,-9483.8,25593.
1324.000000000,5480.5,2321.4,-9481.7,25593.
1325.000000000,5480.6,2321.4,-9480.2,25593.
1326.000000000,5480.6,2321.4,-9478.3,25593.
1327.000000000,5480.7,2321.5,-9476.1,25593.
1328.000000000,5480.8,2321.5,-9476.9,25594.
1329.000000000,5480.8,2321.5,-9476.2,25594.
1330.000000000,5480.9,2321.5,-9475.0,25594.
1331.000000000,5481.0,2321.5,-9473.7,25594.
1332.000000000,5481.0,2321.6,-9471.6,25594.
1333.000000000,5481.1,2321.6,-9469.2,25594.
1334.000000000,5481.2,2321.6,-9466.7,25594.
1335.000000000,5481.2,2321.6,-9464.0,25595.
1336.000000000,5481.3,2321.7,-9461.3,25595.
1337.000000000,5481.4,2321.7,-9458.8,25595.
1338.000000000,5481.4,2321.7,-9456.3,25595.
1339.000000000,5481.5,2321.7,-9453.9,25595.
1340.000000000,5481.5,2321.7,-9451.4,25595.
1341.000000000,5481.6,2321.8,-9448.9,25595.
1342.000000000,5481.7,2321.8,-9446.8,25596.
1343.000000000,5481.7,2321.8,-9444.3,25596.
1344.000000000,5481.8,2321.8,-9441.6,25596.
1345.000000000,5481.9,2321.9,-9438.9,25596.
1346.000000000,5481.9,2321.9,-9436.2,25596.
1347.000000000,5482.0,2321.9,-9433.4,25596.
1348.000000000,5482.1,2321.9,-9430.7,25596.
1349.000000000,5482.1,2321.9,-9427.9,25597.
1350.000000000,5482.2,2322.0,-9425.3,25597.
1351.000000000,5482.3,2322.0,-9422.7,25597.
1352.000000000,5482.3,2322.0,-9420.4,25597.
1353.000000000,5482.4,2322.0,-9417.9,25597.
1354.000000000,5482.4,2322.1,-9415.4,25597.
1355.000000000,5482.5,2322.1,-9412.8,25597.
1356.000000000,5482.6,2322.1,-9410.1,25598.
1357.000000000,5482.6,2322.1,-9407.4,25598.
1358.000000000,5482.7,2322.1,-9404.6,25598.
1359.000000000,5482.8,2322.2,-9401.9,25598.
1360.000000000,5482.8,2322.2,-9399.1,25598.
1361.000000000,5482.9,2322.2,-9396.3,25598.
1362.000000000,5483.0,2322.2,-9393.6,25598.
1363.000000000,5483.0,2322.3,-9390.8,25599.
1364.000000000,5483.1,2322.3,-9390.2,25599.
1365.000000000,5483.2,2322.3,-9393.3,25599.
1366.000000000,5483.2,2322.3,-9393.7,25599.
1367.000000000,5483.3,2322.3,-9392.4,25599.
1368.000000000,5483.3,2322.4,-9390.3,25599.
1369.000000000,5483.4,2322.4,-9387.8,25600.
1370.000000000,5483.5,2322.4,-9385.3,25600.
1371.000000000,5483.5,2322.4,-9382.6,25600.
1372.000000000,5483.6,2322.5,-9379.9,25600.
1373.000000000,5483.7,2322.5,-9377.2,25600.
1374.000000000,5483.7,2322.5,-9374.5,25600.
1375.000000000,5483.8,2322.5,-9371.8,25600.
1376.000000000,5483.9,2322.5,-9369.0,25601.
1377.000000000,5483.9,2322.6,-9366.3,25601.
1378.000000000,5484.0,2322.6,-9363.6,25601.
1379.000000000,5484.1,2322.6,-9360.9,25601.
1380.000000000,5484.1,2322.6,-9358.2,25601.
1381.000000000,5484.2,2322.7,-9355.4,25601.
1382.000000000,5484.2,2322.7,-9352.7,25601.
1383.000000000,5484.3,2322.7,-9350.0,25602.
1384.000000000,5484.4,2322.7,-9347.3,25602.
1385.000000000,5484.4,2322.7,-9344.5,25602.
1386.000000000,5484.5,2322.8,-9341.8,25602.
1387.000000000,5484.6,2322.8,-9339.1,25602.
1388.000000000,5484.6,2322.8,-9336.4,25602.
1389.000000000,5484.7,2322.8,-9333.6,25602.
1390.000000000,5484.8,2322.9,-9330.9,25603.
1391.000000000,5484.8,2322.9,-9328.2,25603.
1392.000000000,5484.9,2322.9,-9325.5,25603.
1393.000000000,5485.0,2322.9,-9322.8,25603.
1394.000000000,5485.0,2322.9,-9320.0,25603.
1395.000000000,5485.1,2323.0,-9317.3,25603.
1396.000000000,5485.1,2323.0,-9314.6,25604.
1397.000000000,5485.2,2323.0,-9311.9,25604.
1398.000000000,5485.3,2323.0,-9309.2,25604.
1399.000000000,5485.3,2323.1,-9306.5,25604.
1400.000000000,5485.4,2323.1,-9303.8,25604.
1401.000000000,5485.5,2323.1,-9301.1,25604.
1402.000000000,5485.5,2323.1,-9298.4,25604.
1403.000000000,5485.6,2323.1,-9295.7,25605.
1404.000000000,5485.7,2323.2,-9293.9,25605.
1405.000000000,5485.7,2323.2,-9291.7,25605.
1406.000000000,5485.8,2323.2,-9289.2,25605.
1407.000000000,5485.8,2323.2,-9286.7,25605.
1408.000000000,5485.9,2323.3,-9284.1,25605.
1409.000000000,5486.0,2323.3,-9281.5,25605.
1410.000000000,5486.0,2323.3,-9280.2,25606.
1411.000000000,5486.1,2323.3,-9278.2,25606.
1412.000000000,5486.2,2323.3,-9275.8,25606.
1413.000000000,5486.2,2323.4,-9273.3,25606.
1414.000000000,5486.3,2323.4,-9270.6,25606.
1415.000000000,5486.4,2323.4,-9268.0,25606.
1416.000000000,5486.4,2323.4,-9265.3,25606.
1417.000000000,5486.5,2323.5,-9262.7,25607.
1418.000000000,5486.6,2323.5,-9260.0,25607.
1419.000000000,5486.6,2323.5,-9257.3,25607.
1420.000000000,5486.7,2323.5,-9254.6,25607.
1421.000000000,5486.7,2323.5,-9252.0,25607.
1422.000000000,5486.8,2323.6,-9249.3,25607.
1423.000000000,5486.9,2323.6,-9246.6,25607.
1424.000000000,5486.9,2323.6,-9243.9,25608.
1425.000000000,5487.0,2323.6,-9241.3,25608.
1426.000000000,5487.1,2323.7,-9238.7,25608.
1427.000000000,5487.1,2323.7,-9236.1,25608.
1428.000000000,5487.2,2323.7,-9233.5,25608.
1429.000000000,5487.3,2323.7,-9230.8,25608.
1430.000000000,5487.3,2323.7,-9228.2,25608.
1431.000000000,5487.4,2323.8,-9225.5,25609.
1432.000000000,5487.5,2323.8,-9222.9,25609.
1433.000000000,5487.5,2323.8,-9220.8,25609.
1434.000000000,5487.6,2323.8,-9219.3,25609.
1435.000000000,5487.6,2323.9,-9220.2,25609.
1436.000000000,5487.7,2323.9,-9219.5,25609.
1437.000000000,5487.8,2323.9,-9217.6,25609.
1438.000000000,5487.8,2323.9,-9215.4,25610.
1439.000000000,5487.9,2324.0,-9212.9,25610.
1440.000000000,5488.0,2324.0,-9210.3,25610.
1441.000000000,5488.0,2324.0,-9207.7,25610.
1442.000000000,5488.1,2324.0,-9205.1,25610.
1443.000000000,5488.2,2324.0,-9202.6,25610.
1444.000000000,5488.2,2324.1,-9200.0,25610.
1445.000000000,5488.3,2324.1,-9197.3,25611.
1446.000000000,5488.4,2324.1,-9194.7,25611.
1447.000000000,5488.4,2324.1,-9192.1,25611.
1448.000000000,5488.5,2324.2,-9189.5,25611.
1449.000000000,5488.5,2324.2,-9186.8,25611.
1450.000000000,5488.6,2324.2,-9184.2,25611.
1451.000000000,5488.7,2324.2,-9181.6,25612.
1452.000000000,5488.7,2324.2,-9179.0,25612.
1453.000000000,5488.8,2324.3,-9176.4,25612.
1454.000000000,5488.9,2324.3,-9173.9,25612.
1455.000000000,5488.9,2324.3,-9171.3,25612.
1456.000000000,5489.0,2324.3,-9168.7,25612.
1457.000000000,5489.1,2324.4,-9166.1,25612.
1458.000000000,5489.1,2324.4,-9163.4,25613.
1459.000000000,5489.2,2324.4,-9160.8,25613.
1460.000000000,5489.3,2324.4,-9158.2,25613.
1461.000000000,5489.3,2324.4,-9155.6,25613.
1462.000000000,5489.4,2324.5,-9152.9,25613.
1463.000000000,5489.5,2324.5,-9150.4,25613.
1464.000000000,5489.5,2324.5,-9147.8,25613.
1465.000000000,5489.6,2324.5,-9145.2,25614.
1466.000000000,5489.6,2324.6,-9142.6,25614.
1467.000000000,5489.7,2324.6,-9140.0,25614.
1468.000000000,5489.8,2324.6,-9137.3,25614.
1469.000000000,5489.8,2324.6,-9134.7,25614.
1470.000000000,5489.9,2324.7,-9132.1,25614.
1471.000000000,5490.0,2324.7,-9129.5,25614.
1472.000000000,5490.0,2324.7,-9126.8,25615.
1473.000000000,5490.1,2324.7,-9124.2,25615.
1474.000000000,5490.2,2324.7,-9121.6,25615.
1475.000000000,5490.2,2324.8,-9119.1,25615.
1476.000000000,5490.3,2324.8,-9116.8,25615.
1477.000000000,5490.4,2324.8,-9114.8,25615.
1478.000000000,5490.4,2324.8,-9112.5,25615.
1479.000000000,5490.5,2324.9,-9110.6,25616.
1480.000000000,5490.6,2324.9,-9108.4,25616.
1481.000000000,5490.6,2324.9,-9105.9,25616.
1482.000000000,5490.7,2324.9,-9103.4,25616.
1483.000000000,5490.8,2324.9,-9100.8,25616.
1484.000000000,5490.8,2325.0,-9098.2,25616.
1485.000000000,5490.9,2325.0,-9095.6,25616.
1486.000000000,5491.0,2325.0,-9093.0,25617.
1487.000000000,5491.0,2325.0,-9090.4,25617.
1488.000000000,5491.1,2325.1,-9087.8,25617.
1489.000000000,5491.1,2325.1,-9085.3,25617.
1490.000000000,5491.2,2325.1,-9082.7,25617.
1491.000000000,5491.3,2325.1,-9080.1,25617.
1492.000000000,5491.3,2325.2,-9077.5,25618.
1493.000000000,5491.4,2325.2,-9074.9,25618.
1494.000000000,5491.5,2325.2,-9072.3,25618.
1495.000000000,5491.5,2325.2,-9069.7,25618.
1496.000000000,5491.6,2325.2,-9067.2,25618.
1497.000000000,5491.7,2325.3,-9064.6,25618.
1498.000000000,5491.7,2325.3,-9062.0,25618.
1499.000000000,5491.8,2325.3,-9059.4,25619.
1500.000000000,5491.9,2325.3,-9056.9,25619.
1501.000000000,5491.9,2325.4,-9054.3,25619.
1502.000000000,5492.0,2325.4,-9051.7,25619.
1503.000000000,5492.1,2325.4,-9049.1,25619.
1504.000000000,5492.1,2325.4,-9046.5,25619.
1505.000000000,5492.2,2325.5,-9044.0,25619.
1506.000000000,5492.3,2325.5,-9043.5,25620.
1507.000000000,5492.3,2325.5,-9041.9,25620.
1508.000000000,5492.4,2325.5,-9039.7,25620.
1509.000000000,5492.5,2325.5,-9037.3,25620.
1510.000000000,5492.5,2325.6,-9034.9,25620.
1511.000000000,5492.6,2325.6,-9032.4,25620.
1512.000000000,5492.7,2325.6,-9030.1,25620.
1513.000000000,5492.7,2325.6,-9027.7,25621.
1514.000000000,5492.8,2325.7,-9025.2,25621.
1515.000000000,5492.8,2325.7,-9022.7,25621.
1516.000000000,5492.9,2325.7,-9020.2,25621.
1517.000000000,5493.0,2325.7,-9017.6,25621.
1518.000000000,5493.0,2325.8,-9015.1,25621.
1519.000000000,5493.1,2325.8,-9012.5,25621.
1520.000000000,5493.2,2325.8,-9010.0,25622.
1521.000000000,5493.2,2325.8,-9007.4,25622.
1522.000000000,5493.3,2325.8,-9004.9,25622.
1523.000000000,5493.4,2325.9,-9002.4,25622.
1524.000000000,5493.4,2325.9,-8999.8,25622.
1525.000000000,5493.5,2325.9,-8997.4,25622.
1526.000000000,5493.6,2325.9,-8995.0,25622.
1527.000000000,5493.6,2326.0,-8992.5,25623.
1528.000000000,5493.7,2326.0,-8990.0,25623.
1529.000000000,5493.8,2326.0,-8987.4,25623.
1530.000000000,5493.8,2326.0,-8984.9,25623.
1531.000000000,5493.9,2326.1,-8982.4,25623.
1532.000000000,5494.0,2326.1,-8979.9,25623.
1533.000000000,5494.0,2326.1,-8977.4,25624.
1534.000000000,5494.1,2326.1,-8974.9,25624.
1535.000000000,5494.2,2326.1,-8972.4,25624.
1536.000000000,5494.2,2326.2,-8969.8,25624.
1537.000000000,5494.3,2326.2,-8967.3,25624.
1538.000000000,5494.4,2326.2,-8964.8,25624.
1539.000000000,5494.4,2326.2,-8962.3,25624.
1540.000000000,5494.5,2326.3,-8959.8,25625.
1541.000000000,5494.6,2326.3,-8957.2,25625.
1542.000000000,5494.6,2326.3,-8954.7,25625.
1543.000000000,5494.7,2326.3,-8952.2,25625.
1544.000000000,5494.8,2326.4,-8949.7,25625.
1545.000000000,5494.8,2326.4,-8947.2,25625.
1546.000000000,5494.9,2326.4,-8944.7,25625.
1547.000000000,5495.0,2326.4,-8942.2,25626.
1548.000000000,5495.0,2326.4,-8939.7,25626.
1549.000000000,5495.1,2326.5,-8938.2,25626.
1550.000000000,5495.2,2326.5,-8936.1,25626.
1551.000000000,5495.2,2326.5,-8933.7,25626.
1552.000000000,5495.3,2326.5,-8931.3,25626.
1553.000000000,5495.4,2326.6,-8930.7,25626.
1554.000000000,5495.4,2326.6,-8929.0,25627.
1555.000000000,5495.5,2326.6,-8926.8,25627.
1556.000000000,5495.6,2326.6,-8924.5,25627.
1557.000000000,5495.6,2326.7,-8922.1,25627.
1558.000000000,5495.7,2326.7,-8919.6,25627.
1559.000000000,5495.8,2326.7,-8917.2,25627.
1560.000000000,5495.8,2326.7,-8914.7,25627.
1561.000000000,5495.9,2326.7,-8912.2,25628.
1562.000000000,5495.9,2326.8,-8910.3,25628.
1563.000000000,5496.0,2326.8,-8908.2,25628.
1564.000000000,5496.1,2326.8,-8906.1,25628.
1565.000000000,5496.1,2326.8,-8904.6,25628.
1566.000000000,5496.2,2326.9,-8902.6,25628.
1567.000000000,5496.3,2326.9,-8900.3,25628.
1568.000000000,5496.3,2326.9,-8898.3,25629.
1569.000000000,5496.4,2326.9,-8896.0,25629.
1570.000000000,5496.5,2327.0,-8893.6,25629.
1571.000000000,5496.5,2327.0,-8891.1,25629.
1572.000000000,5496.6,2327.0,-8888.7,25629.
1573.000000000,5496.7,2327.0,-8886.2,25629.
1574.000000000,5496.7,2327.1,-8883.8,25629.
1575.000000000,5496.8,2327.1,-8881.3,25630.
1576.000000000,5496.9,2327.1,-8878.9,25630.
1577.000000000,5496.9,2327.1,-8876.4,25630.
1578.000000000,5497.0,2327.1,-8874.0,25630.
1579.000000000,5497.1,2327.2,-8871.5,25630.
1580.000000000,5497.1,2327.2,-8869.1,25630.
1581.000000000,5497.2,2327.2,-8866.6,25630.
1582.000000000,5497.3,2327.2,-8864.2,25631.
1583.000000000,5497.3,2327.3,-8861.7,25631.
1584.000000000,5497.4,2327.3,-8859.3,25631.
1585.000000000,5497.5,2327.3,-8856.8,25631.
1586.000000000,5497.5,2327.3,-8854.4,25631.
1587.000000000,5497.6,2327.4,-8851.9,25631.
1588.000000000,5497.7,2327.4,-8849.5,25631.
1589.000000000,5497.7,2327.4,-8847.1,25632.
1590.000000000,5497.8,2327.4,-8844.6,25632.
1591.000000000,5497.9,2327.4,-8842.2,25632.
1592.000000000,5497.9,2327.5,-8840.5,25632.
1593.000000000,5498.0,2327.5,-8838.4,25632.
1594.000000000,5498.1,2327.5,-8836.1,25632.
1595.000000000,5498.1,2327.5,-8833.7,25632.
1596.000000000,5498.2,2327.6,-8831.3,25633.
1597.000000000,5498.3,2327.6,-8828.9,25633.
1598.000000000,5498.3,2327.6,-8826.5,25633.
1599.000000000,5498.4,2327.6,-8824.1,25633.
1600.000000000,5498.5,2327.7,-8821.7,25633.
1601.000000000,5498.5,2327.7,-8820.7,25633.
1602.000000000,5498.6,2327.7,-8819.0,25634.
1603.000000000,5498.7,2327.7,-8818.1,25634.
1604.000000000,5498.7,2327.8,-8816.4,25634.
1605.000000000,5498.8,2327.8,-8814.3,25634.
1606.000000000,5498.9,2327.8,-8812.1,25634.
1607.000000000,5498.9,2327.8,-8809.7,25634.
1608.000000000,5499.0,2327.8,-8807.4,25634.
1609.000000000,5499.1,2327.9,-8805.0,25635.
1610.000000000,5499.1,2327.9,-8804.0,25635.
1611.000000000,5499.2,2327.9,-8802.3,25635.
1612.000000000,5499.3,2327.9,-8804.9,25635.
1613.000000000,5499.3,2328.0,-8805.3,25635.
1614.000000000,5499.4,2328.0,-8804.3,25635.
1615.000000000,5499.5,2328.0,-8802.8,25635.
1616.000000000,5499.5,2328.0,-8801.7,25636.
1617.000000000,5499.6,2328.1,-8800.0,25636.
1618.000000000,5499.7,2328.1,-8797.9,25636.
1619.000000000,5499.7,2328.1,-8795.7,25636.
1620.000000000,5499.8,2328.1,-8793.4,25636.
1621.000000000,5499.9,2328.2,-8791.0,25636.
1622.000000000,5499.9,2328.2,-8788.7,25636.
1623.000000000,5500.0,2328.2,-8786.3,25636.
1624.000000000,5500.1,2328.2,-8784.0,25637.
1625.000000000,5500.1,2328.2,-8781.6,25637.
1626.000000000,5500.2,2328.3,-8779.2,25637.
1627.000000000,5500.3,2328.3,-8776.8,25637.
1628.000000000,5500.3,2328.3,-8774.5,25637.
1629.000000000,5500.4,2328.3,-8772.1,25637.
1630.000000000,5500.5,2328.4,-8769.7,25638.
1631.000000000,5500.5,2328.4,-8767.3,25638.
1632.000000000,5500.6,2328.4,-8765.0,25638.
1633.000000000,5500.7,2328.4,-8762.6,25638.
1634.000000000,5500.7,2328.5,-8760.2,25638.
1635.000000000,5500.8,2328.5,-8757.8,25638.
1636.000000000,5500.9,2328.5,-8755.5,25638.
1637.000000000,5500.9,2328.5,-8753.1,25639.
1638.000000000,5501.0,2328.6,-8750.8,25639.
1639.000000000,5501.1,2328.6,-8748.8,25639.
1640.000000000,5501.1,2328.6,-8746.7,25639.
1641.000000000,5501.2,2328.6,-8744.4,25639.
1642.000000000,5501.3,2328.6,-8742.1,25639.
1643.000000000,5501.3,2328.7,-8739.8,25639.
1644.000000000,5501.4,2328.7,-8737.4,25640.
1645.000000000,5501.5,2328.7,-8735.1,25640.
1646.000000000,5501.5,2328.7,-8732.7,25640.
1647.000000000,5501.6,2328.8,-8730.4,25640.
1648.000000000,5501.7,2328.8,-8728.1,25640.
1649.000000000,5501.7,2328.8,-8726.4,25640.
1650.000000000,5501.8,2328.8,-8725.0,25640.
1651.000000000,5501.9,2328.9,-8723.0,25641.
1652.000000000,5501.9,2328.9,-8720.8,25641.
1653.000000000,5502.0,2328.9,-8718.6,25641.
1654.000000000,5502.1,2328.9,-8716.2,25641.
1655.000000000,5502.1,2329.0,-8713.9,25641.
1656.000000000,5502.2,2329.0,-8711.7,25641.
1657.000000000,5502.3,2329.0,-8709.7,25641.
1658.000000000,5502.3,2329.0,-8707.8,25642.
1659.000000000,5502.4,2329.1,-8705.9,25642.
1660.000000000,5502.5,2329.1,-8703.8,25642.
1661.000000000,5502.5,2329.1,-8701.7,25642.
1662.000000000,5502.6,2329.1,-8699.4,25642.
1663.000000000,5502.7,2329.1,-8697.1,25642.
1664.000000000,5502.7,2329.2,-8694.8,25642.
1665.000000000,5502.8,2329.2,-8692.4,25643.
1666.000000000,5502.9,2329.2,-8691.5,25643.
1667.000000000,5502.9,2329.2,-8689.8,25643.
1668.000000000,5503.0,2329.3,-8687.7,25643.
1669.000000000,5503.1,2329.3,-8685.5,25643.
1670.000000000,5503.1,2329.3,-8683.2,25643.
1671.000000000,5503.2,2329.3,-8680.9,25643.
1672.000000000,5503.3,2329.4,-8678.6,25644.
1673.000000000,5503.3,2329.4,-8676.4,25644.
1674.000000000,5503.4,2329.4,-8674.2,25644.
1675.000000000,5503.5,2329.4,-8672.2,25644.
1676.000000000,5503.5,2329.5,-8670.3,25644.
1677.000000000,5503.6,2329.5,-8668.1,25644.
1678.000000000,5503.7,2329.5,-8665.9,25644.
1679.000000000,5503.7,2329.5,-8663.6,25645.
1680.000000000,5503.8,2329.6,-8661.3,25645.
1681.000000000,5503.9,2329.6,-8659.1,25645.
1682.000000000,5503.9,2329.6,-8658.6,25645.
1683.000000000,5504.0,2329.6,-8657.1,25645.
1684.000000000,5504.1,2329.6,-8655.1,25645.
1685.000000000,5504.1,2329.7,-8653.0,25645.
1686.000000000,5504.2,2329.7,-8650.7,25646.
1687.000000000,5504.3,2329.7,-8648.5,25646.
1688.000000000,5504.3,2329.7,-8646.2,25646.
1689.000000000,5504.4,2329.8,-8644.0,25646.
1690.000000000,5504.5,2329.8,-8641.8,25646.
1691.000000000,5504.5,2329.8,-8639.5,25646.
1692.000000000,5504.6,2329.8,-8637.2,25646.
1693.000000000,5504.7,2329.9,-8634.9,25647.
1694.000000000,5504.7,2329.9,-8632.6,25647.
1695.000000000,5504.8,2329.9,-8630.3,25647.
1696.000000000,5504.9,2329.9,-8628.0,25647.
1697.000000000,5504.9,2330.0,-8626.1,25647.
1698.000000000,5505.0,2330.0,-8624.6,25647.
1699.000000000,5505.1,2330.0,-8622.6,25647.
1700.000000000,5505.1,2330.0,-8620.8,25648.
1701.000000000,5505.2,2330.1,-8618.8,25648.
1702.000000000,5505.3,2330.1,-8616.6,25648.
1703.000000000,5505.3,2330.1,-8614.3,25648.
1704.000000000,5505.4,2330.1,-8612.0,25648.
1705.000000000,5505.5,2330.2,-8609.7,25648.
1706.000000000,5505.5,2330.2,-8607.4,25648.
1707.000000000,5505.6,2330.2,-8605.2,25649.
1708.000000000,5505.7,2330.2,-8602.9,25649.
1709.000000000,5505.7,2330.2,-8600.6,25649.
1710.000000000,5505.8,2330.3,-8598.3,25649.
1711.000000000,5505.9,2330.3,-8596.0,25649.
1712.000000000,5505.9,2330.3,-8593.7,25649.
1713.000000000,5506.0,2330.3,-8591.4,25649.
1714.000000000,5506.1,2330.4,-8589.1,25650.
1715.000000000,5506.2,2330.4,-8586.9,25650.
1716.000000000,5506.2,2330.4,-8584.6,25650.
1717.000000000,5506.3,2330.4,-8582.3,25650.
1718.000000000,5506.4,2330.5,-8580.0,25650.
1719.000000000,5506.4,2330.5,-8577.7,25650.
1720.000000000,5506.5,2330.5,-8575.4,25650.
1721.000000000,5506.6,2330.5,-8573.1,25651.
1722.000000000,5506.6,2330.6,-8570.9,25651.
1723.000000000,5506.7,2330.6,-8568.6,25651.
1724.000000000,5506.8,2330.6,-8566.3,25651.
1725.000000000,5506.8,2330.6,-8564.1,25651.
1726.000000000,5506.9,2330.7,-8561.8,25651.
1727.000000000,5507.0,2330.7,-8559.6,25651.
1728.000000000,5507.0,2330.7,-8557.3,25652.
1729.000000000,5507.1,2330.7,-8556.6,25652.
1730.000000000,5507.2,2330.8,-8556.0,25652.
1731.000000000,5507.2,2330.8,-8557.6,25652.
1732.000000000,5507.3,2330.8,-8560.1,25652.
1733.000000000,5507.4,2330.8,-8561.3,25652.
1734.000000000,5507.4,2330.9,-8561.1,25652.
1735.000000000,5507.5,2330.9,-8559.9,25653.
1736.000000000,5507.6,2330.9,-8558.1,25653.
1737.000000000,5507.6,2330.9,-8556.1,25653.
1738.000000000,5507.7,2330.9,-8554.9,25653.
1739.000000000,5507.8,2331.0,-8553.3,25653.
1740.000000000,5507.8,2331.0,-8551.3,25653.
1741.000000000,5507.9,2331.0,-8549.2,25653.
1742.000000000,5508.0,2331.0,-8547.0,25654.
1743.000000000,5508.0,2331.1,-8544.8,25654.
1744.000000000,5508.1,2331.1,-8543.1,25654.
1745.000000000,5508.2,2331.1,-8541.1,25654.
1746.000000000,5508.2,2331.1,-8539.0,25654.
1747.000000000,5508.3,2331.2,-8536.8,25654.
1748.000000000,5508.4,2331.2,-8534.6,25654.
1749.000000000,5508.4,2331.2,-8532.4,25655.
1750.000000000,5508.5,2331.2,-8530.2,25655.
1751.000000000,5508.6,2331.3,-8527.9,25655.
1752.000000000,5508.6,2331.3,-8525.7,25655.
1753.000000000,5508.7,2331.3,-8523.5,25655.
1754.000000000,5508.8,2331.3,-8521.2,25655.
1755.000000000,5508.8,2331.4,-8519.0,25655.
1756.000000000,5508.9,2331.4,-8516.8,25656.
1757.000000000,5509.0,2331.4,-8514.5,25656.
1758.000000000,5509.0,2331.4,-8512.3,25656.
1759.000000000,5509.1,2331.5,-8510.0,25656.
1760.000000000,5509.2,2331.5,-8507.8,25656.
1761.000000000,5509.2,2331.5,-8505.6,25656.
1762.000000000,5509.3,2331.5,-8503.3,25656.
1763.000000000,5509.4,2331.6,-8501.1,25656.
1764.000000000,5509.4,2331.6,-8498.9,25657.
1765.000000000,5509.5,2331.6,-8496.6,25657.
1766.000000000,5509.6,2331.6,-8494.4,25657.
1767.000000000,5509.6,2331.7,-8492.2,25657.
1768.000000000,5509.7,2331.7,-8490.0,25657.
1769.000000000,5509.8,2331.7,-8487.7,25657.
1770.000000000,5509.8,2331.7,-8485.5,25657.
1771.000000000,5509.9,2331.8,-8483.3,25658.
1772.000000000,5510.0,2331.8,-8481.0,25658.
1773.000000000,5510.0,2331.8,-8478.8,25658.
1774.000000000,5510.1,2331.8,-8476.6,25658.
1775.000000000,5510.2,2331.8,-8474.4,25658.
1776.000000000,5510.2,2331.9,-8472.2,25658.
1777.000000000,5510.3,2331.9,-8470.1,25658.
1778.000000000,5510.4,2331.9,-8467.9,25659.
1779.000000000,5510.4,2331.9,-8465.8,25659.
1780.000000000,5510.5,2332.0,-8463.6,25659.
1781.000000000,5510.6,2332.0,-8461.4,25659.
1782.000000000,5510.6,2332.0,-8459.2,25659.
1783.000000000,5510.7,2332.0,-8457.0,25659.
1784.000000000,5510.8,2332.1,-8454.8,25659.
1785.000000000,5510.8,2332.1,-8452.6,25660.
1786.000000000,5510.9,2332.1,-8450.3,25660.
1787.000000000,5510.9,2332.1,-8448.1,25660.
1788.000000000,5511.0,2332.2,-8445.9,25660.
1789.000000000,5511.1,2332.2,-8443.7,25660.
1790.000000000,5511.1,2332.2,-8441.5,25660.
1791.000000000,5511.2,2332.2,-8439.3,25660.
1792.000000000,5511.3,2332.3,-8437.1,25661.
1793.000000000,5511.3,2332.3,-8434.9,25661.
1794.000000000,5511.4,2332.3,-8432.7,25661.
1795.000000000,5511.5,2332.3,-8430.5,25661.
1796.000000000,5511.5,2332.4,-8428.2,25661.
1797.000000000,5511.6,2332.4,-8426.0,25661.
1798.000000000,5511.7,2332.4,-8423.8,25661.
1799.000000000,5511.7,2332.4,-8421.6,25662.
1800.000000000,5511.8,2332.5,-8419.4,25662.
1801.000000000,5511.9,2332.5,-8417.7,25662.
1802.000000000,5511.9,2332.5,-8417.2,25662.
1803.000000000,5512.0,2332.5,-8416.2,25662.
1804.000000000,5512.1,2332.6,-8414.5,25662.
1805.000000000,5512.1,2332.6,-8412.6,25662.
1806.000000000,5512.2,2332.6,-8410.5,25663.
1807.000000000,5512.3,2332.6,-8408.3,25663.
1808.000000000,5512.3,2332.7,-8406.2,25663.
1809.000000000,5512.4,2332.7,-8404.0,25663.
1810.000000000,5512.4,2332.7,-8401.8,25663.
1811.000000000,5512.5,2332.7,-8399.7,25663.
1812.000000000,5512.6,2332.8,-8398.1,25663.
1813.000000000,5512.6,2332.8,-8396.2,25664.
1814.000000000,5512.7,2332.8,-8394.2,25664.
1815.000000000,5512.8,2332.8,-8392.1,25664.
1816.000000000,5512.8,2332.9,-8390.0,25664.
1817.000000000,5512.9,2332.9,-8387.9,25664.
1818.000000000,5513.0,2332.9,-8385.7,25664.
1819.000000000,5513.0,2332.9,-8383.6,25664.
1820.000000000,5513.1,2332.9,-8381.4,25664.
1821.000000000,5513.2,2333.0,-8379.3,25665.
1822.000000000,5513.2,2333.0,-8377.2,25665.
1823.000000000,5513.3,2333.0,-8375.1,25665.
1824.000000000,5513.4,2333.0,-8372.9,25665.
1825.000000000,5513.4,2333.1,-8370.8,25665.
1826.000000000,5513.5,2333.1,-8368.6,25665.
1827.000000000,5513.6,2333.1,-8366.5,25665.
1828.000000000,5513.6,2333.1,-8364.4,25666.
1829.000000000,5513.7,2333.2,-8362.2,25666.
1830.000000000,5513.8,2333.2,-8360.1,25666.
1831.000000000,5513.8,2333.2,-8357.9,25666.
1832.000000000,5513.9,2333.2,-8355.8,25666.
1833.000000000,5514.0,2333.3,-8353.6,25666.
1834.000000000,5514.0,2333.3,-8351.5,25666.
1835.000000000,5514.1,2333.3,-8349.3,25667.
1836.000000000,5514.1,2333.3,-8347.2,25667.
1837.000000000,5514.2,2333.4,-8345.1,25667.
1838.000000000,5514.3,2333.4,-8342.9,25667.
1839.000000000,5514.3,2333.4,-8340.8,25667.
1840.000000000,5514.4,2333.4,-8338.7,25667.
1841.000000000,5514.5,2333.5,-8336.5,25667.
1842.000000000,5514.5,2333.5,-8334.4,25668.
1843.000000000,5514.6,2333.5,-8332.3,25668.
1844.000000000,5514.7,2333.5,-8330.2,25668.
1845.000000000,5514.7,2333.6,-8328.1,25668.
1846.000000000,5514.8,2333.6,-8326.0,25668.
1847.000000000,5514.9,2333.6,-8323.9,25668.
1848.000000000,5514.9,2333.6,-8321.8,25668.
1849.000000000,5515.0,2333.7,-8319.7,25669.
1850.000000000,5515.1,2333.7,-8317.5,25669.
1851.000000000,5515.1,2333.7,-8315.4,25669.
1852.000000000,5515.2,2333.7,-8313.3,25669.
1853.000000000,5515.3,2333.8,-8311.2,25669.
1854.000000000,5515.3,2333.8,-8309.1,25669.
1855.000000000,5515.4,2333.8,-8307.0,25669.
1856.000000000,5515.5,2333.8,-8304.8,25670.
1857.000000000,5515.5,2333.9,-8302.7,25670.
1858.000000000,5515.6,2333.9,-8300.6,25670.
1859.000000000,5515.7,2333.9,-8298.5,25670.
1860.000000000,5515.7,2333.9,-8296.4,25670.
1861.000000000,5515.8,2334.0,-8294.3,25670.
1862.000000000,5515.9,2334.0,-8292.2,25670.
1863.000000000,5515.9,2334.0,-8290.1,25670.
1864.000000000,5516.0,2334.0,-8288.1,25671.
1865.000000000,5516.1,2334.1,-8286.0,25671.
1866.000000000,5516.1,2334.1,-8283.9,25671.
1867.000000000,5516.2,2334.1,-8281.8,25671.
1868.000000000,5516.3,2334.1,-8279.7,25671.
1869.000000000,5516.3,2334.2,-8277.6,25671.
1870.000000000,5516.4,2334.2,-8275.6,25671.
1871.000000000,5516.4,2334.2,-8273.6,25672.
1872.000000000,5516.5,2334.2,-8271.5,25672.
1873.000000000,5516.6,2334.3,-8269.4,25672.
1874.000000000,5516.6,2334.3,-8267.3,25672.
1875.000000000,5516.7,2334.3,-8265.2,25672.
1876.000000000,5516.8,2334.3,-8263.3,25672.
1877.000000000,5516.8,2334.4,-8261.7,25672.
1878.000000000,5516.9,2334.4,-8261.7,25673.
1879.000000000,5517.0,2334.4,-8260.6,25673.
1880.000000000,5517.0,2334.4,-8259.0,25673.
1881.000000000,5517.1,2334.5,-8257.1,25673.
1882.000000000,5517.2,2334.5,-8255.2,25673.
1883.000000000,5517.2,2334.5,-8253.2,25673.
1884.000000000,5517.3,2334.5,-8251.1,25673.
1885.000000000,5517.4,2334.6,-8249.1,25674.
1886.000000000,5517.4,2334.6,-8247.1,25674.
1887.000000000,5517.5,2334.6,-8245.1,25674.
1888.000000000,5517.6,2334.6,-8243.0,25674.
1889.000000000,5517.6,2334.7,-8241.0,25674.
1890.000000000,5517.7,2334.7,-8238.9,25674.
1891.000000000,5517.8,2334.7,-8236.8,25674.
1892.000000000,5517.8,2334.7,-8234.8,25675.
1893.000000000,5517.9,2334.8,-8232.7,25675.
1894.000000000,5518.0,2334.8,-8230.6,25675.
1895.000000000,5518.0,2334.8,-8228.6,25675.
1896.000000000,5518.1,2334.8,-8226.5,25675.
1897.000000000,5518.2,2334.9,-8224.5,25675.
1898.000000000,5518.2,2334.9,-8222.4,25675.
1899.000000000,5518.3,2334.9,-8220.3,25676.
1900.000000000,5518.4,2334.9,-8218.3,25676.
1901.000000000,5518.4,2335.0,-8216.2,25676.
1902.000000000,5518.5,2335.0,-8214.2,25676.
1903.000000000,5518.6,2335.0,-8212.1,25676.
1904.000000000,5518.6,2335.0,-8210.1,25676.
1905.000000000,5518.7,2335.1,-8208.0,25676.
1906.000000000,5518.8,2335.1,-8206.0,25676.
1907.000000000,5518.8,2335.1,-8203.9,25677.
1908.000000000,5518.9,2335.1,-8201.9,25677.
1909.000000000,5519.0,2335.2,-8199.8,25677.
1910.000000000,5519.0,2335.2,-8197.8,25677.
1911.000000000,5519.1,2335.2,-8195.7,25677.
1912.000000000,5519.2,2335.2,-8193.7,25677.
1913.000000000,5519.2,2335.3,-8191.7,25677.
1914.000000000,5519.3,2335.3,-8189.7,25678.
1915.000000000,5519.4,2335.3,-8187.7,25678.
1916.000000000,5519.4,2335.3,-8185.6,25678.
1917.000000000,5519.5,2335.4,-8183.6,25678.
1918.000000000,5519.6,2335.4,-8181.6,25678.
1919.000000000,5519.6,2335.4,-8179.5,25678.
1920.000000000,5519.7,2335.4,-8177.5,25678.
1921.000000000,5519.8,2335.5,-8175.4,25679.
1922.000000000,5519.8,2335.5,-8173.4,25679.
1923.000000000,5519.9,2335.5,-8171.4,25679.
1924.000000000,5520.0,2335.5,-8169.3,25679.
1925.000000000,5520.0,2335.6,-8167.3,25679.
1926.000000000,5520.1,2335.6,-8165.3,25679.
1927.000000000,5520.2,2335.6,-8163.3,25679.
1928.000000000,5520.2,2335.6,-8161.2,25680.
1929.000000000,5520.3,2335.7,-8159.2,25680.
1930.000000000,5520.4,2335.7,-8157.2,25680.
1931.000000000,5520.4,2335.7,-8155.2,25680.
1932.000000000,5520.5,2335.7,-8153.2,25680.
1933.000000000,5520.6,2335.8,-8151.2,25680.
1934.000000000,5520.6,2335.8,-8149.2,25680.
1935.000000000,5520.7,2335.8,-8147.2,25681.
1936.000000000,5520.8,2335.8,-8145.2,25681.
1937.000000000,5520.8,2335.9,-8143.2,25681.
1938.000000000,5520.9,2335.9,-8141.2,25681.
1939.000000000,5521.0,2335.9,-8139.2,25681.
1940.000000000,5521.0,2335.9,-8137.2,25681.
1941.000000000,5521.1,2336.0,-8135.2,25681.
1942.000000000,5521.2,2336.0,-8133.4,25681.
1943.000000000,5521.2,2336.0,-8131.6,25682.
1944.000000000,5521.3,2336.0,-8129.6,25682.
1945.000000000,5521.4,2336.1,-8127.6,25682.
1946.000000000,5521.4,2336.1,-8125.7,25682.
1947.000000000,5521.5,2336.1,-8123.7,25682.
1948.000000000,5521.6,2336.1,-8121.7,25682.
1949.000000000,5521.6,2336.2,-8119.8,25682.
1950.000000000,5521.7,2336.2,-8119.9,25683.
1951.000000000,5521.8,2336.2,-8119.1,25683.
1952.000000000,5521.8,2336.2,-8117.7,25683.
1953.000000000,5521.9,2336.3,-8116.0,25683.
1954.000000000,5522.0,2336.3,-8114.1,25683.
1955.000000000,5522.0,2336.3,-8112.2,25683.
1956.000000000,5522.1,2336.3,-8110.2,25683.
1957.000000000,5522.2,2336.4,-8108.3,25684.
1958.000000000,5522.2,2336.4,-8106.3,25684.
1959.000000000,5522.3,2336.4,-8104.3,25684.
1960.000000000,5522.4,2336.4,-8102.3,25684.
1961.000000000,5522.4,2336.5,-8100.3,25684.
1962.000000000,5522.5,2336.5,-8098.4,25684.
1963.000000000,5522.6,2336.5,-8096.4,25684.
1964.000000000,5522.7,2336.5,-8094.4,25685.
1965.000000000,5522.7,2336.6,-8092.4,25685.
1966.000000000,5522.8,2336.6,-8090.7,25685.
1967.000000000,5522.9,2336.6,-8090.7,25685.
1968.000000000,5522.9,2336.6,-8089.7,25685.
1969.000000000,5523.0,2336.7,-8088.2,25685.
1970.000000000,5523.1,2336.7,-8086.4,25685.
1971.000000000,5523.1,2336.7,-8084.5,25685.
1972.000000000,5523.2,2336.7,-8082.6,25686.
1973.000000000,5523.3,2336.8,-8080.6,25686.
1974.000000000,5523.3,2336.8,-8078.7,25686.
1975.000000000,5523.4,2336.8,-8076.7,25686.
1976.000000000,5523.5,2336.8,-8074.7,25686.
1977.000000000,5523.5,2336.9,-8072.8,25686.
1978.000000000,5523.6,2336.9,-8070.8,25686.
1979.000000000,5523.7,2336.9,-8068.8,25687.
1980.000000000,5523.7,2337.0,-8066.9,25687.
1981.000000000,5523.8,2337.0,-8065.0,25687.
1982.000000000,5523.9,2337.0,-8063.1,25687.
1983.000000000,5523.9,2337.0,-8061.2,25687.
1984.000000000,5524.0,2337.1,-8059.2,25687.
1985.000000000,5524.1,2337.1,-8057.2,25687.
1986.000000000,5524.1,2337.1,-8055.3,25688.
1987.000000000,5524.2,2337.1,-8053.3,25688.
1988.000000000,5524.3,2337.2,-8051.4,25688.
1989.000000000,5524.3,2337.2,-8049.4,25688.
1990.000000000,5524.4,2337.2,-8047.5,25688.
1991.000000000,5524.5,2337.2,-8045.5,25688.
1992.000000000,5524.5,2337.3,-8043.5,25688.
1993.000000000,5524.6,2337.3,-8041.6,25689.
1994.000000000,5524.7,2337.3,-8039.6,25689.
1995.000000000,5524.8,2337.3,-8037.7,25689.
1996.000000000,5524.8,2337.4,-8035.9,25689.
1997.000000000,5524.9,2337.4,-8034.0,25689.
1998.000000000,5525.0,2337.4,-8032.1,25689.
1999.000000000,5525.0,2337.4,-8030.2,25689.
2000.000000000,5525.1,2337.5,-8028.2,25689.
2001.000000000,5525.2,2337.5,-8026.3,25690.
2002.000000000,5525.2,2337.5,-8024.4,25690.
2003.000000000,5525.3,2337.5,-8022.4,25690.
2004.000000000,5525.4,2337.6,-8020.5,25690.
2005.000000000,5525.4,2337.6,-8018.5,25690.
2006.000000000,5525.5,2337.6,-8016.6,25690.
2007.000000000,5525.6,2337.6,-8014.8,25690.
2008.000000000,5525.6,2337.7,-8012.9,25691.
2009.000000000,5525.7,2337.7,-8011.0,25691.
2010.000000000,5525.8,2337.7,-8009.0,25691.
2011.000000000,5525.8,2337.7,-8007.1,25691.
2012.000000000,5525.9,2337.8,-8005.4,25691.
2013.000000000,5526.0,2337.8,-8003.9,25691.
2014.000000000,5526.0,2337.8,-8003.0,25691.
2015.000000000,5526.1,2337.8,-8002.4,25692.
2016.000000000,5526.2,2337.9,-8001.5,25692.
2017.000000000,5526.3,2337.9,-8000.6,25692.
2018.000000000,5526.3,2337.9,-7999.2,25692.
2019.000000000,5526.4,2337.9,-7997.5,25692.
2020.000000000,5526.5,2338.0,-7995.6,25692.
2021.000000000,5526.5,2338.0,-7993.8,25692.
2022.000000000,5526.6,2338.0,-7991.9,25693.
2023.000000000,5526.7,2338.0,-7990.0,25693.
2024.000000000,5526.7,2338.1,-7988.1,25693.
2025.000000000,5526.8,2338.1,-7986.1,25693.
2026.000000000,5526.9,2338.1,-7984.2,25693.
2027.000000000,5526.9,2338.1,-7982.3,25693.
2028.000000000,5527.0,2338.2,-7980.4,25693.
2029.000000000,5527.1,2338.2,-7978.5,25694.
2030.000000000,5527.1,2338.2,-7976.6,25694.
2031.000000000,5527.2,2338.3,-7974.7,25694.
2032.000000000,5527.3,2338.3,-7972.7,25694.
2033.000000000,5527.3,2338.3,-7970.8,25694.
2034.000000000,5527.4,2338.3,-7968.9,25694.
2035.000000000,5527.5,2338.4,-7967.0,25694.
2036.000000000,5527.6,2338.4,-7965.1,25694.
2037.000000000,5527.6,2338.4,-7963.2,25695.
2038.000000000,5527.7,2338.4,-7963.3,25695.
2039.000000000,5527.8,2338.5,-7962.4,25695.
2040.000000000,5527.8,2338.5,-7960.9,25695.
2041.000000000,5527.9,2338.5,-7959.2,25695.
2042.000000000,5528.0,2338.5,-7957.4,25695.
2043.000000000,5528.0,2338.6,-7955.5,25695.
2044.000000000,5528.1,2338.6,-7953.6,25696.
2045.000000000,5528.2,2338.6,-7951.7,25696.
2046.000000000,5528.2,2338.6,-7949.8,25696.
2047.000000000,5528.3,2338.7,-7947.9,25696.
2048.000000000,5528.4,2338.7,-7946.1,25696.
2049.000000000,5528.4,2338.7,-7944.9,25696.
2050.000000000,5528.5,2338.7,-7943.9,25696.
2051.000000000,5528.6,2338.8,-7943.1,25697.
2052.000000000,5528.7,2338.8,-7941.9,25697.
2053.000000000,5528.7,2338.8,-7940.3,25697.
2054.000000000,5528.8,2338.8,-7938.5,25697.
2055.000000000,5528.9,2338.9,-7936.7,25697.
2056.000000000,5528.9,2338.9,-7934.9,25697.
2057.000000000,5529.0,2338.9,-7933.0,25697.
2058.000000000,5529.1,2338.9,-7931.3,25698.
2059.000000000,5529.1,2339.0,-7929.8,25698.
2060.000000000,5529.2,2339.0,-7928.1,25698.
2061.000000000,5529.3,2339.0,-7926.3,25698.
2062.000000000,5529.3,2339.0,-7924.5,25698.
2063.000000000,5529.4,2339.1,-7922.6,25698.
2064.000000000,5529.5,2339.1,-7920.8,25698.
2065.000000000,5529.5,2339.1,-7918.9,25698.
2066.000000000,5529.6,2339.2,-7917.0,25699.
2067.000000000,5529.7,2339.2,-7915.1,25699.
2068.000000000,5529.7,2339.2,-7913.3,25699.
2069.000000000,5529.8,2339.2,-7911.4,25699.
